CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 30 100 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 86 325 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 87 263 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
7 Ground~
168 340 172 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
9 Inverter~
13 215 391 0 2 22
0 3 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
6153 0 0
0
0
2 +V
167 454 441 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
14 Logic Display~
6 1016 472 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 931 473 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 961 472 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 989 474 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 898 475 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 813 476 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 843 475 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 871 477 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
7 74LS273
150 559 468 0 18 37
0 6 4 23 22 21 20 19 18 17
16 14 13 12 11 10 9 8 7
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U5
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
7 Ground~
168 708 354 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7668 0 0
0
0
6 74LS83
105 492 364 0 14 29
0 14 13 12 11 27 26 25 24 15
22 21 20 19 23
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
6 74LS83
105 620 366 0 14 29
0 10 9 8 7 2 2 2 2 2
18 17 16 40 15
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U3
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
14 Logic Display~
6 444 91 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
9 2-In AND~
219 596 194 0 3 22
0 36 32 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 1 0
1 U
3789 0 0
0
0
9 2-In AND~
219 656 193 0 3 22
0 35 32 26
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
4871 0 0
0
0
9 2-In AND~
219 713 194 0 3 22
0 34 32 25
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3750 0 0
0
0
9 2-In AND~
219 771 194 0 3 22
0 33 32 24
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
8778 0 0
0
0
6 74LS95
110 387 116 0 12 25
0 5 3 3 31 30 29 28 2 32
39 38 37
0
0 0 13040 0
6 74LS95
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
538 0 0
0
0
14 Logic Display~
6 585 37 0 1 2
10 36
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 615 36 0 1 2
10 35
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
14 Logic Display~
6 643 38 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5950 0 0
0
0
14 Logic Display~
6 670 36 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 304 48 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 277 50 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6735 0 0
0
0
14 Logic Display~
6 249 48 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8365 0 0
0
0
14 Logic Display~
6 219 49 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4132 0 0
0
0
10 Ascii Key~
169 819 126 0 11 12
0 33 34 35 36 41 42 43 44 0
0 53
0
0 0 4656 602
0
4 KBD2
-12 -39 16 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 0 0 0 0
3 KBD
4551 0 0
0
0
10 Ascii Key~
169 118 169 0 11 12
0 31 30 29 28 45 46 47 48 0
0 55
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 0 0 0 0
3 KBD
3635 0 0
0
0
62
8 1 2 0 0 4096 0 23 3 0 0 3
355 152
340 152
340 166
1 0 3 0 0 8192 0 4 0 0 5 3
200 391
174 391
174 325
2 2 4 0 0 12416 0 4 14 0 0 5
236 391
346 391
346 421
527 421
527 441
3 0 3 0 0 0 0 23 0 0 5 2
349 107
327 107
1 2 3 0 0 4224 0 1 23 0 0 4
98 325
327 325
327 98
349 98
1 1 5 0 0 4224 0 23 2 0 0 4
355 89
164 89
164 263
99 263
1 1 6 0 0 8320 0 14 5 0 0 6
518 435
518 425
446 425
446 458
454 458
454 450
0 1 7 0 0 4224 0 0 6 22 0 3
599 539
1016 539
1016 490
1 0 8 0 0 8320 0 9 0 0 23 3
989 492
989 529
590 529
0 1 9 0 0 4224 0 0 8 24 0 3
581 518
961 518
961 490
1 0 10 0 0 8320 0 7 0 0 25 3
931 491
931 511
572 511
1 0 11 0 0 8320 0 10 0 0 26 4
898 493
898 614
526 614
526 529
1 0 12 0 0 8320 0 13 0 0 27 4
871 495
871 605
516 605
516 520
0 1 13 0 0 8320 0 0 12 28 0 4
507 513
507 597
843 597
843 493
0 1 14 0 0 8320 0 0 11 29 0 4
500 505
500 588
813 588
813 494
9 0 2 0 0 4096 0 17 0 0 20 2
663 336
663 311
8 0 2 0 0 0 0 17 0 0 20 2
645 336
645 311
7 0 2 0 0 0 0 17 0 0 20 2
636 336
636 311
6 0 2 0 0 0 0 17 0 0 20 2
627 336
627 311
1 5 2 0 0 8320 0 15 17 0 0 4
708 348
708 311
618 311
618 336
14 9 15 0 0 8320 0 17 16 0 0 5
663 400
663 428
549 428
549 334
535 334
4 18 7 0 0 0 0 17 14 0 0 6
609 336
609 275
372 275
372 571
599 571
599 505
17 3 8 0 0 0 0 14 17 0 0 6
590 505
590 559
379 559
379 284
600 284
600 336
2 16 9 0 0 0 0 17 14 0 0 6
591 336
591 292
387 292
387 550
581 550
581 505
15 1 10 0 0 0 0 14 17 0 0 6
572 505
572 539
396 539
396 301
582 301
582 336
4 14 11 0 0 0 0 16 14 0 0 6
481 334
481 309
406 309
406 529
563 529
563 505
13 3 12 0 0 0 0 14 16 0 0 6
554 505
554 520
415 520
415 317
472 317
472 334
2 12 13 0 0 0 0 16 14 0 0 6
463 334
463 325
424 325
424 513
545 513
545 505
11 1 14 0 0 0 0 14 16 0 0 4
536 505
431 505
431 334
454 334
12 10 16 0 0 8320 0 17 14 0 0 4
627 400
627 420
599 420
599 441
11 9 17 0 0 12416 0 17 14 0 0 4
618 400
618 411
590 411
590 441
8 10 18 0 0 4224 0 14 17 0 0 4
581 441
581 405
609 405
609 400
13 7 19 0 0 8320 0 16 14 0 0 4
508 398
508 404
572 404
572 441
12 6 20 0 0 8320 0 16 14 0 0 4
499 398
499 408
563 408
563 441
11 5 21 0 0 8320 0 16 14 0 0 4
490 398
490 413
554 413
554 441
10 4 22 0 0 8320 0 16 14 0 0 4
481 398
481 417
545 417
545 441
14 3 23 0 0 8320 0 16 14 0 0 3
535 398
536 398
536 441
3 8 24 0 0 8320 0 22 16 0 0 4
769 217
769 235
517 235
517 334
3 7 25 0 0 8320 0 21 16 0 0 4
711 217
711 229
508 229
508 334
3 6 26 0 0 8320 0 20 16 0 0 4
654 216
654 223
499 223
499 334
3 5 27 0 0 8320 0 19 16 0 0 3
594 217
490 217
490 334
7 0 28 0 0 4224 0 23 0 0 49 2
355 143
219 143
6 0 29 0 0 4224 0 23 0 0 48 2
355 134
249 134
5 0 30 0 0 4096 0 23 0 0 45 2
355 125
277 125
1 2 30 0 0 8320 0 29 33 0 0 3
277 68
277 153
143 153
4 0 31 0 0 8192 0 23 0 0 47 3
355 116
355 117
304 117
1 1 31 0 0 4224 0 33 28 0 0 3
143 147
304 147
304 66
3 1 29 0 0 0 0 33 30 0 0 3
143 159
249 159
249 66
4 1 28 0 0 0 0 33 31 0 0 3
143 165
219 165
219 67
2 0 32 0 0 4096 0 19 0 0 53 2
585 172
585 151
2 0 32 0 0 0 0 20 0 0 53 2
645 171
645 151
2 0 32 0 0 0 0 21 0 0 53 2
702 172
702 151
9 2 32 0 0 12416 0 23 22 0 0 5
419 125
561 125
561 151
760 151
760 172
1 0 33 0 0 4096 0 22 0 0 62 2
778 172
778 104
1 0 34 0 0 4096 0 21 0 0 61 2
720 172
720 110
1 0 35 0 0 4096 0 20 0 0 60 2
663 171
663 116
1 0 36 0 0 4096 0 19 0 0 59 2
603 172
603 122
1 9 32 0 0 128 0 18 23 0 0 3
444 109
444 125
419 125
4 1 36 0 0 4224 0 32 24 0 0 3
794 122
585 122
585 55
3 1 35 0 0 4224 0 32 25 0 0 3
794 116
615 116
615 54
2 1 34 0 0 4224 0 32 26 0 0 3
794 110
643 110
643 56
1 1 33 0 0 8320 0 27 32 0 0 3
670 54
670 104
794 104
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
