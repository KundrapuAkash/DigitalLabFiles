CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
19
14 Logic Display~
6 530 260 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 496 258 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 461 259 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 565 259 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 918 134 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 1025 137 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 991 135 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 956 136 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 1060 136 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
7 Ground~
168 716 304 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7931 0 0
0
0
6 74LS83
105 768 228 0 14 29
0 12 13 14 15 8 9 10 11 2
3 4 5 6 7
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
14 Logic Display~
6 565 115 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 496 114 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 461 115 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 530 116 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
2 +V
167 268 306 0 1 3
0 20
0
0 0 54256 180
2 5V
7 -2 21 6
2 V1
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4718 0 0
0
0
7 Buffer~
58 213 250 0 2 22
0 22 21
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3874 0 0
0
0
7 74LS273
150 319 221 0 18 37
0 20 21 12 13 14 15 16 17 18
19 8 9 10 11 12 13 14 15
0
0 0 13040 692
7 74LS273
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
10 Ascii Key~
169 137 230 0 11 12
0 19 18 17 16 23 24 25 22 0
0 57
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 0 0 0 0
3 KBD
3789 0 0
0
0
33
10 1 3 0 0 4224 0 11 8 0 0 3
800 219
956 219
956 154
11 1 4 0 0 4224 0 11 7 0 0 3
800 228
991 228
991 153
12 1 5 0 0 4224 0 11 6 0 0 3
800 237
1025 237
1025 155
13 1 6 0 0 4224 0 11 9 0 0 3
800 246
1060 246
1060 154
14 1 7 0 0 8320 0 11 5 0 0 3
800 273
918 273
918 152
9 1 2 0 0 8320 0 11 10 0 0 3
736 273
716 273
716 298
0 5 8 0 0 8320 0 0 11 18 0 5
451 288
451 346
630 346
630 228
736 228
0 6 9 0 0 16512 0 0 11 17 0 5
488 298
488 333
603 333
603 237
736 237
0 7 10 0 0 12288 0 0 11 16 0 4
530 301
594 301
594 246
736 246
8 0 11 0 0 4096 0 11 0 0 15 4
736 255
587 255
587 293
565 293
0 1 12 0 0 4224 0 0 11 23 0 5
461 207
618 207
618 185
736 185
736 192
0 2 13 0 0 8320 0 0 11 24 0 3
495 198
495 201
736 201
0 3 14 0 0 4096 0 0 11 25 0 4
530 189
653 189
653 210
736 210
0 4 15 0 0 12288 0 0 11 26 0 4
565 180
642 180
642 219
736 219
14 1 11 0 0 12416 0 18 4 0 0 5
351 216
388 216
388 322
565 322
565 277
13 1 10 0 0 12416 0 18 1 0 0 5
351 225
377 225
377 308
530 308
530 278
12 1 9 0 0 128 0 18 2 0 0 5
351 234
364 234
364 298
496 298
496 276
11 1 8 0 0 128 0 18 3 0 0 4
351 243
351 288
461 288
461 277
0 3 12 0 0 128 0 0 18 23 0 5
378 207
378 118
243 118
243 243
287 243
0 4 13 0 0 0 0 0 18 24 0 5
370 198
370 129
253 129
253 234
287 234
0 5 14 0 0 0 0 0 18 25 0 5
361 189
361 139
263 139
263 225
287 225
18 6 15 0 0 0 0 18 18 0 0 5
351 180
351 152
273 152
273 216
287 216
15 1 12 0 0 128 0 18 14 0 0 3
351 207
461 207
461 133
16 1 13 0 0 128 0 18 13 0 0 3
351 198
496 198
496 132
17 1 14 0 0 4224 0 18 15 0 0 3
351 189
530 189
530 134
18 1 15 0 0 4224 0 18 12 0 0 3
351 180
565 180
565 133
4 7 16 0 0 12416 0 19 18 0 0 4
162 226
195 226
195 207
287 207
3 8 17 0 0 12416 0 19 18 0 0 4
162 220
185 220
185 198
287 198
2 9 18 0 0 12416 0 19 18 0 0 4
162 214
173 214
173 189
287 189
1 10 19 0 0 8320 0 19 18 0 0 3
162 208
162 180
287 180
1 1 20 0 0 8320 0 18 16 0 0 3
281 261
268 261
268 291
2 2 21 0 0 4224 0 17 18 0 0 4
228 250
273 250
273 252
287 252
8 1 22 0 0 4224 0 19 17 0 0 2
162 250
198 250
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
