CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 29 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
31
7 Ground~
168 280 394 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
6 74LS90
107 266 341 0 10 21
0 2 56 2 57 5 4 58 59 60
4
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U9
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
4441 0 0
0
0
7 Ground~
168 229 273 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 252 69 0 1 3
0 7
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
9 CA 7-Seg~
184 253 169 0 18 19
10 2 2 4 61 2 2 2 62 6
0 0 2 2 0 0 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5394 0 0
0
0
7 Ground~
168 500 392 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
2 +V
167 459 75 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
9 CA 7-Seg~
184 459 163 0 18 19
10 19 18 17 16 13 14 15 63 20
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3747 0 0
0
0
6 74LS90
107 479 344 0 10 21
0 2 64 5 8 9 5 11 12 10
5
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U8
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
6 74LS47
187 444 256 0 14 29
0 11 12 10 5 65 66 15 14 13
16 17 18 19 67
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U7
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
7 Ground~
168 646 393 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
6 74LS47
187 590 256 0 14 29
0 9 23 8 22 68 69 26 25 24
27 28 29 30 70
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U5
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
6 74LS90
107 626 338 0 10 21
0 2 71 5 8 21 22 9 23 8
22
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U6
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
9 CA 7-Seg~
184 605 163 0 18 19
10 30 29 28 27 24 25 26 72 31
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3363 0 0
0
0
2 +V
167 605 75 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
7 Ground~
168 770 409 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
2 +V
167 720 74 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
9 CA 7-Seg~
184 720 162 0 18 19
10 43 42 41 40 37 38 39 73 44
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6671 0 0
0
0
6 74LS90
107 743 336 0 10 21
0 2 74 21 32 33 35 36 21 32
35
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U4
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
0
0
6 74LS47
187 705 255 0 14 29
0 36 21 32 35 75 76 39 38 37
40 41 42 43 77
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U3
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4871 0 0
0
0
6 74LS47
187 834 252 0 14 29
0 33 46 47 45 78 79 50 49 48
51 52 53 54 80
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
6 74LS90
107 872 333 0 10 21
0 2 81 2 82 34 45 33 46 47
45
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U2
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
8778 0 0
0
0
9 CA 7-Seg~
184 849 159 0 18 19
10 54 53 52 51 48 49 50 83 55
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
538 0 0
0
0
2 +V
167 849 71 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6843 0 0
0
0
7 Ground~
168 906 378 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3136 0 0
0
0
7 Pulser~
4 821 445 0 10 12
0 84 85 34 86 0 0 5 5 6
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5950 0 0
0
0
9 Resistor~
219 253 103 0 4 5
0 6 7 0 1
0
0 0 880 90
3 150
7 0 28 8
2 R5
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 459 105 0 4 5
0 20 3 0 1
0
0 0 880 90
3 150
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 605 105 0 4 5
0 31 3 0 1
0
0 0 880 90
3 150
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 720 104 0 4 5
0 44 3 0 1
0
0 0 880 90
3 150
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 849 101 0 4 5
0 55 3 0 1
0
0 0 880 90
3 150
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
83
3 0 4 0 0 4224 0 5 0 0 5 3
244 205
244 295
227 295
5 0 5 0 0 8192 0 2 0 0 15 3
242 373
242 418
410 418
3 1 2 0 0 4096 0 2 1 0 0 3
269 367
269 388
280 388
1 1 2 0 0 0 0 2 1 0 0 3
287 367
287 388
280 388
6 10 4 0 0 0 0 2 2 0 0 6
233 373
233 377
219 377
219 295
233 295
233 303
7 0 2 0 0 4096 0 5 0 0 7 3
268 205
268 253
262 253
6 0 2 0 0 4096 0 5 0 0 8 3
262 205
262 258
256 258
5 0 2 0 0 4096 0 5 0 0 9 3
256 205
256 260
238 260
2 0 2 0 0 4096 0 5 0 0 10 3
238 205
238 263
232 263
1 1 2 0 0 4224 0 5 3 0 0 3
232 205
232 267
229 267
1 9 6 0 0 4224 0 27 5 0 0 2
253 121
253 133
1 2 7 0 0 8320 0 4 27 0 0 3
252 78
253 78
253 85
4 0 8 0 0 8320 0 9 0 0 14 4
473 370
473 429
606 429
606 383
9 4 8 0 0 0 0 13 13 0 0 5
611 300
606 300
606 383
620 383
620 364
3 0 5 0 0 8320 0 13 0 0 16 4
629 364
629 506
410 506
410 396
0 3 5 0 0 0 0 0 9 20 0 5
428 343
397 343
397 396
482 396
482 370
7 5 9 0 0 12416 0 13 9 0 0 5
647 300
667 300
667 473
455 473
455 376
1 1 2 0 0 0 0 9 6 0 0 2
500 370
500 386
3 9 10 0 0 4224 0 10 9 0 0 3
467 293
467 306
464 306
6 10 5 0 0 0 0 9 9 0 0 4
446 376
428 376
428 306
446 306
1 7 11 0 0 8320 0 10 9 0 0 4
485 293
485 291
500 291
500 306
2 8 12 0 0 4224 0 10 9 0 0 3
476 293
476 306
482 306
4 10 5 0 0 0 0 10 9 0 0 4
458 293
458 299
446 299
446 306
5 9 13 0 0 12416 0 8 10 0 0 4
462 199
462 205
467 205
467 223
6 8 14 0 0 12416 0 8 10 0 0 4
468 199
468 205
476 205
476 223
7 7 15 0 0 12416 0 8 10 0 0 4
474 199
474 202
485 202
485 223
4 10 16 0 0 12416 0 8 10 0 0 4
456 199
456 205
458 205
458 223
3 11 17 0 0 12416 0 8 10 0 0 4
450 199
450 203
449 203
449 223
2 12 18 0 0 12416 0 8 10 0 0 4
444 199
444 203
440 203
440 223
1 13 19 0 0 12416 0 8 10 0 0 4
438 199
438 203
431 203
431 223
1 9 20 0 0 4224 0 28 8 0 0 2
459 123
459 127
1 2 3 0 0 4224 0 7 28 0 0 2
459 84
459 87
5 0 21 0 0 8320 0 13 0 0 51 4
602 370
602 412
751 412
751 385
3 9 8 0 0 0 0 12 13 0 0 3
613 293
613 300
611 300
6 10 22 0 0 8320 0 13 13 0 0 4
593 370
574 370
574 300
593 300
1 1 2 0 0 0 0 13 11 0 0 5
647 364
647 381
644 381
644 387
646 387
1 7 9 0 0 0 0 12 13 0 0 4
631 293
631 291
647 291
647 300
2 8 23 0 0 4224 0 12 13 0 0 3
622 293
622 300
629 300
4 10 22 0 0 0 0 12 13 0 0 4
604 293
604 299
593 299
593 300
5 9 24 0 0 12416 0 14 12 0 0 4
608 199
608 205
613 205
613 223
6 8 25 0 0 12416 0 14 12 0 0 4
614 199
614 205
622 205
622 223
7 7 26 0 0 12416 0 14 12 0 0 4
620 199
620 202
631 202
631 223
4 10 27 0 0 12416 0 14 12 0 0 4
602 199
602 205
604 205
604 223
3 11 28 0 0 12416 0 14 12 0 0 4
596 199
596 203
595 203
595 223
2 12 29 0 0 12416 0 14 12 0 0 4
590 199
590 203
586 203
586 223
1 13 30 0 0 12416 0 14 12 0 0 4
584 199
584 203
577 203
577 223
1 9 31 0 0 4224 0 29 14 0 0 2
605 123
605 127
1 2 3 0 0 0 0 15 29 0 0 2
605 84
605 87
1 1 2 0 0 0 0 19 16 0 0 4
764 362
764 395
770 395
770 403
4 9 32 0 0 12416 0 19 19 0 0 5
737 362
737 389
672 389
672 298
728 298
3 8 21 0 0 0 0 19 19 0 0 6
746 362
746 385
794 385
794 295
746 295
746 298
7 5 33 0 0 12416 0 22 19 0 0 4
893 295
918 295
918 368
719 368
5 3 34 0 0 4224 0 22 26 0 0 5
848 365
848 423
859 423
859 436
845 436
6 10 35 0 0 12416 0 19 19 0 0 6
710 368
710 372
696 372
696 290
710 290
710 298
1 7 36 0 0 8320 0 20 19 0 0 4
746 292
746 287
764 287
764 298
2 8 21 0 0 0 0 20 19 0 0 4
737 292
737 287
746 287
746 298
3 9 32 0 0 0 0 20 19 0 0 4
728 292
728 287
728 287
728 298
4 10 35 0 0 0 0 20 19 0 0 4
719 292
719 287
710 287
710 298
5 9 37 0 0 12416 0 18 20 0 0 4
723 198
723 204
728 204
728 222
6 8 38 0 0 12416 0 18 20 0 0 4
729 198
729 204
737 204
737 222
7 7 39 0 0 12416 0 18 20 0 0 4
735 198
735 201
746 201
746 222
4 10 40 0 0 12416 0 18 20 0 0 4
717 198
717 204
719 204
719 222
3 11 41 0 0 12416 0 18 20 0 0 4
711 198
711 202
710 202
710 222
2 12 42 0 0 12416 0 18 20 0 0 4
705 198
705 202
701 202
701 222
1 13 43 0 0 12416 0 18 20 0 0 4
699 198
699 202
692 202
692 222
1 9 44 0 0 4224 0 30 18 0 0 2
720 122
720 126
1 2 3 0 0 0 0 17 30 0 0 2
720 83
720 86
6 10 45 0 0 12416 0 22 22 0 0 6
839 365
839 369
825 369
825 287
839 287
839 295
3 1 2 0 0 0 0 22 25 0 0 3
875 359
875 372
906 372
1 1 2 0 0 0 0 22 25 0 0 3
893 359
893 372
906 372
1 7 33 0 0 0 0 21 22 0 0 4
875 289
875 288
893 288
893 295
2 8 46 0 0 8320 0 21 22 0 0 4
866 289
866 297
875 297
875 295
3 9 47 0 0 12416 0 21 22 0 0 4
857 289
857 284
857 284
857 295
4 10 45 0 0 0 0 21 22 0 0 4
848 289
848 297
839 297
839 295
5 9 48 0 0 12416 0 23 21 0 0 4
852 195
852 201
857 201
857 219
6 8 49 0 0 12416 0 23 21 0 0 4
858 195
858 201
866 201
866 219
7 7 50 0 0 12416 0 23 21 0 0 4
864 195
864 198
875 198
875 219
4 10 51 0 0 12416 0 23 21 0 0 4
846 195
846 201
848 201
848 219
3 11 52 0 0 12416 0 23 21 0 0 4
840 195
840 199
839 199
839 219
2 12 53 0 0 12416 0 23 21 0 0 4
834 195
834 199
830 199
830 219
1 13 54 0 0 12416 0 23 21 0 0 4
828 195
828 199
821 199
821 219
1 9 55 0 0 4224 0 31 23 0 0 2
849 119
849 123
1 2 3 0 0 0 0 24 31 0 0 2
849 80
849 83
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
