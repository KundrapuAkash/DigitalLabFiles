CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
23
8 2-In OR~
219 840 249 0 3 22
0 6 5 8
0
0 0 624 512
6 74LS32
-21 -24 21 -16
3 U6B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
8953 0 0
0
0
8 2-In OR~
219 730 251 0 3 22
0 4 9 3
0
0 0 624 512
6 74LS32
-21 -24 21 -16
3 U6A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 161454668
65 0 0 0 4 1 3 0
1 U
4441 0 0
0
0
9 Inverter~
13 671 315 0 2 22
0 3 10
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U8A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
3618 0 0
0
0
6 74LS47
187 396 401 0 14 29
0 11 12 13 14 38 39 21 20 19
18 17 16 15 40
0
0 0 13040 512
6 74LS47
-21 -60 21 -52
2 U7
-2 -61 12 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6153 0 0
0
0
9 CA 7-Seg~
184 219 314 0 18 19
10 41 10 10 42 43 44 45 46 22
2 1 1 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5394 0 0
0
0
9 CA 7-Seg~
184 310 314 0 18 19
10 15 16 17 18 19 20 21 47 22
2 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7734 0 0
0
0
9 2-In AND~
219 784 259 0 3 22
0 8 7 9
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1348791995
65 0 0 0 4 1 2 0
1 U
9914 0 0
0
0
7 Ground~
168 769 425 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
6 74LS83
105 853 378 0 14 29
0 7 5 6 23 2 3 3 2 2
11 12 13 14 48
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
7 Ground~
168 609 259 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
14 Logic Display~
6 361 131 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 395 130 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 430 130 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 464 129 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 460 34 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 426 35 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 391 35 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 357 36 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
2 +V
167 220 199 0 1 3
0 22
0
0 0 54256 180
2 5V
7 -2 21 6
2 V1
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
10 Ascii Key~
169 124 97 0 11 12
0 37 36 35 34 49 50 51 33 0
0 48
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
4871 0 0
0
0
7 Buffer~
58 203 149 0 2 22
0 33 32
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3750 0 0
0
0
7 74LS273
150 263 118 0 18 37
0 22 32 28 29 30 31 34 35 36
37 27 26 25 24 28 29 30 31
0
0 0 13040 692
7 74LS273
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
6 74LS83
105 650 190 0 14 29
0 28 29 30 31 27 26 25 24 2
7 5 6 23 4
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
538 0 0
0
0
59
1 0 3 0 0 8192 0 3 0 0 24 3
692 315
692 316
703 316
6 0 3 0 0 4096 0 9 0 0 24 3
846 348
846 316
837 316
14 1 4 0 0 8320 0 23 2 0 0 5
682 235
682 216
753 216
753 242
749 242
2 0 5 0 0 4096 0 1 0 0 29 2
859 258
882 258
1 0 6 0 0 4096 0 1 0 0 30 4
859 240
877 240
877 239
873 239
2 0 7 0 0 4096 0 7 0 0 28 2
804 268
891 268
1 3 8 0 0 8320 0 7 1 0 0 3
804 250
804 249
813 249
2 3 9 0 0 8320 0 2 7 0 0 3
749 260
749 259
759 259
3 0 10 0 0 4096 0 5 0 0 10 3
210 350
210 379
204 379
2 2 10 0 0 8320 0 3 5 0 0 4
656 315
656 509
204 509
204 350
10 1 11 0 0 8320 0 9 4 0 0 5
864 412
864 480
488 480
488 365
434 365
11 2 12 0 0 8320 0 9 4 0 0 5
855 412
855 472
497 472
497 374
434 374
12 3 13 0 0 8320 0 9 4 0 0 5
846 412
846 461
507 461
507 383
434 383
13 4 14 0 0 8320 0 9 4 0 0 5
837 412
837 453
514 453
514 392
434 392
1 13 15 0 0 8320 0 6 4 0 0 3
289 350
289 419
364 419
2 12 16 0 0 8320 0 6 4 0 0 3
295 350
295 410
364 410
3 11 17 0 0 8320 0 6 4 0 0 3
301 350
301 401
364 401
4 10 18 0 0 8320 0 6 4 0 0 3
307 350
307 392
364 392
5 9 19 0 0 8320 0 6 4 0 0 3
313 350
313 383
364 383
6 8 20 0 0 8320 0 6 4 0 0 3
319 350
319 374
364 374
7 7 21 0 0 8320 0 6 4 0 0 3
325 350
325 365
364 365
0 9 22 0 0 4224 0 0 6 23 0 3
207 245
310 245
310 278
1 9 22 0 0 0 0 19 5 0 0 5
220 184
207 184
207 273
219 273
219 278
7 3 3 0 0 8320 0 9 2 0 0 4
837 348
837 316
703 316
703 251
9 0 2 0 0 4096 0 9 0 0 27 2
810 348
810 329
5 0 2 0 0 8192 0 9 0 0 27 3
855 348
855 329
828 329
8 1 2 0 0 12416 0 9 8 0 0 4
828 348
828 329
769 329
769 419
10 1 7 0 0 4224 0 23 9 0 0 3
682 181
891 181
891 348
2 11 5 0 0 8320 0 9 23 0 0 3
882 348
882 190
682 190
12 3 6 0 0 4224 0 23 9 0 0 3
682 199
873 199
873 348
13 4 23 0 0 4224 0 23 9 0 0 3
682 208
864 208
864 348
9 1 2 0 0 0 0 23 10 0 0 3
618 235
609 235
609 253
1 0 24 0 0 4096 0 14 0 0 40 2
464 147
464 217
1 0 25 0 0 4096 0 13 0 0 39 2
430 148
430 208
1 0 26 0 0 4096 0 12 0 0 38 2
395 148
395 199
1 0 27 0 0 4096 0 11 0 0 37 2
361 149
361 190
5 11 27 0 0 4224 0 23 22 0 0 3
618 190
295 190
295 140
12 6 26 0 0 12416 0 22 23 0 0 4
295 131
308 131
308 199
618 199
7 13 25 0 0 4224 0 23 22 0 0 4
618 208
316 208
316 122
295 122
8 14 24 0 0 4224 0 23 22 0 0 4
618 217
323 217
323 113
295 113
1 0 28 0 0 4096 0 18 0 0 45 2
357 54
357 104
1 0 29 0 0 4096 0 17 0 0 46 2
391 53
391 95
1 0 30 0 0 4096 0 16 0 0 47 2
426 53
426 86
1 0 31 0 0 4096 0 15 0 0 48 2
460 52
460 77
15 1 28 0 0 4224 0 22 23 0 0 4
295 104
585 104
585 154
618 154
16 2 29 0 0 4224 0 22 23 0 0 4
295 95
577 95
577 163
618 163
17 3 30 0 0 4224 0 22 23 0 0 4
295 86
570 86
570 172
618 172
18 4 31 0 0 4224 0 22 23 0 0 4
295 77
563 77
563 181
618 181
17 5 30 0 0 0 0 22 22 0 0 6
295 86
303 86
303 31
206 31
206 122
231 122
4 16 29 0 0 0 0 22 22 0 0 6
231 131
219 131
219 20
310 20
310 95
295 95
3 15 28 0 0 0 0 22 22 0 0 6
231 140
223 140
223 15
317 15
317 104
295 104
18 6 31 0 0 0 0 22 22 0 0 5
295 77
295 49
212 49
212 113
231 113
1 1 22 0 0 0 0 22 19 0 0 3
225 158
220 158
220 184
2 2 32 0 0 4224 0 21 22 0 0 2
218 149
231 149
8 1 33 0 0 8320 0 20 21 0 0 4
149 117
180 117
180 149
188 149
4 7 34 0 0 4224 0 20 22 0 0 4
149 93
217 93
217 104
231 104
3 8 35 0 0 4224 0 20 22 0 0 4
149 87
217 87
217 95
231 95
2 9 36 0 0 4224 0 20 22 0 0 4
149 81
217 81
217 86
231 86
1 10 37 0 0 4224 0 20 22 0 0 4
149 75
217 75
217 77
231 77
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
