CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
20
9 Inverter~
13 567 594 0 2 22
0 3 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 1 0
1 U
8953 0 0
0
0
9 Inverter~
13 568 514 0 2 22
0 5 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 1 0
1 U
4441 0 0
0
0
10 3-In NAND~
219 770 555 0 4 22
0 6 7 4 8
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 6 0
1 U
3618 0 0
0
0
2 +V
167 923 58 0 1 3
0 15
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
9 CA 7-Seg~
184 923 133 0 18 19
10 8 9 10 11 12 13 14 28 15
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5394 0 0
0
0
8 3-In OR~
219 591 308 0 4 22
0 21 22 23 26
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 5 0
1 U
7734 0 0
0
0
8 2-In OR~
219 595 122 0 3 22
0 19 20 25
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1580708967
65 0 0 0 4 1 4 0
1 U
9914 0 0
0
0
9 3-In AND~
219 475 86 0 4 22
0 3 7 5 19
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 3 0
1 U
3747 0 0
0
0
9 3-In AND~
219 474 156 0 4 22
0 3 18 16 20
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 3 0
1 U
3549 0 0
0
0
9 3-In AND~
219 474 235 0 4 22
0 17 18 16 21
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
7931 0 0
0
0
9 2-In AND~
219 473 310 0 3 22
0 5 7 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
9325 0 0
0
0
9 2-In AND~
219 474 385 0 3 22
0 7 17 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
8903 0 0
0
0
9 2-In AND~
219 475 464 0 3 22
0 7 16 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1563931748
65 0 0 0 4 1 2 0
1 U
3834 0 0
0
0
9 Inverter~
13 315 359 0 2 22
0 5 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
3363 0 0
0
0
9 Inverter~
13 315 323 0 2 22
0 7 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
7668 0 0
0
0
9 Inverter~
13 316 282 0 2 22
0 3 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
4718 0 0
0
0
6 74LS47
187 774 314 0 14 29
0 23 24 26 25 29 30 14 13 12
11 10 9 8 31
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
7 Ground~
168 165 89 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
6 74LS93
109 232 123 0 8 17
0 2 2 32 27 3 7 5 33
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
0
0
7 Pulser~
4 129 150 0 10 12
0 34 35 27 36 0 0 5 5 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4871 0 0
0
0
44
1 0 3 0 0 8320 0 1 0 0 27 4
552 594
187 594
187 218
289 218
3 2 4 0 0 4224 0 3 1 0 0 3
746 564
588 564
588 594
1 0 5 0 0 4224 0 2 0 0 29 4
553 514
211 514
211 237
272 237
1 2 6 0 0 4224 0 3 2 0 0 4
746 546
592 546
592 514
589 514
2 0 7 0 0 4224 0 3 0 0 28 4
746 555
200 555
200 227
281 227
4 0 8 0 0 8320 0 3 0 0 7 3
797 555
882 555
882 332
13 1 8 0 0 0 0 17 5 0 0 3
812 332
902 332
902 169
12 2 9 0 0 8320 0 17 5 0 0 3
812 323
908 323
908 169
11 3 10 0 0 8320 0 17 5 0 0 3
812 314
914 314
914 169
10 4 11 0 0 8320 0 17 5 0 0 3
812 305
920 305
920 169
9 5 12 0 0 8320 0 17 5 0 0 3
812 296
926 296
926 169
8 6 13 0 0 4224 0 17 5 0 0 3
812 287
932 287
932 169
7 7 14 0 0 4224 0 17 5 0 0 3
812 278
938 278
938 169
1 9 15 0 0 4224 0 4 5 0 0 2
923 67
923 97
2 0 16 0 0 8320 0 13 0 0 22 3
451 473
392 473
392 244
0 2 17 0 0 4224 0 0 12 26 0 3
399 226
399 394
450 394
0 1 7 0 0 0 0 0 12 18 0 3
404 375
404 376
450 376
0 1 7 0 0 0 0 0 13 20 0 3
404 317
404 455
451 455
0 1 5 0 0 0 0 0 11 30 0 3
416 132
416 301
449 301
0 2 7 0 0 0 0 0 11 31 0 3
404 123
404 319
449 319
0 1 3 0 0 0 0 0 9 32 0 3
370 114
370 147
450 147
0 3 16 0 0 0 0 0 9 24 0 3
392 244
392 165
450 165
0 2 18 0 0 4096 0 0 9 25 0 3
381 235
381 156
450 156
2 3 16 0 0 0 0 14 10 0 0 4
336 359
368 359
368 244
450 244
2 2 18 0 0 12416 0 15 10 0 0 4
336 323
356 323
356 235
450 235
2 1 17 0 0 0 0 16 10 0 0 4
337 282
346 282
346 226
450 226
1 0 3 0 0 128 0 16 0 0 32 3
301 282
289 282
289 114
1 0 7 0 0 128 0 15 0 0 31 3
300 323
281 323
281 123
0 1 5 0 0 128 0 0 14 30 0 3
272 132
272 359
300 359
7 3 5 0 0 0 0 19 8 0 0 4
264 132
417 132
417 95
451 95
6 2 7 0 0 0 0 19 8 0 0 4
264 123
407 123
407 86
451 86
5 1 3 0 0 0 0 19 8 0 0 4
264 114
399 114
399 77
451 77
4 1 19 0 0 4224 0 8 7 0 0 4
496 86
574 86
574 113
582 113
4 2 20 0 0 4224 0 9 7 0 0 4
495 156
574 156
574 131
582 131
4 1 21 0 0 4224 0 10 6 0 0 4
495 235
570 235
570 299
578 299
3 2 22 0 0 4224 0 11 6 0 0 4
494 310
570 310
570 308
579 308
0 3 23 0 0 4096 0 0 6 39 0 3
521 385
521 317
578 317
3 2 24 0 0 8320 0 13 17 0 0 4
496 464
668 464
668 287
742 287
3 1 23 0 0 4224 0 12 17 0 0 4
495 385
657 385
657 278
742 278
3 4 25 0 0 8320 0 7 17 0 0 4
628 122
645 122
645 305
742 305
4 3 26 0 0 12416 0 6 17 0 0 4
624 308
636 308
636 296
742 296
1 0 2 0 0 4224 0 19 0 0 43 2
200 114
151 114
2 1 2 0 0 0 0 19 18 0 0 5
200 123
151 123
151 75
165 75
165 83
4 3 27 0 0 4224 0 19 20 0 0 2
194 141
153 141
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
