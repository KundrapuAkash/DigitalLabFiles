CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
39
9 Inverter~
13 962 262 0 2 22
0 3 4
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 6 0
1 U
8953 0 0
0
0
10 2-In NAND~
219 813 206 0 3 22
0 6 8 5
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -642089372
65 0 0 0 4 1 3 0
1 U
4441 0 0
0
0
9 2-In XOR~
219 732 228 0 3 22
0 7 6 8
0
0 0 624 692
6 74LS86
-21 -24 21 -16
4 U10B
-10 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 5 0
1 U
3618 0 0
0
0
8 2-In OR~
219 841 490 0 3 22
0 12 7 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 7 0
1 U
6153 0 0
0
0
9 2-In AND~
219 926 500 0 3 22
0 11 10 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 8 0
1 U
5394 0 0
0
0
9 2-In AND~
219 783 481 0 3 22
0 14 13 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 8 0
1 U
7734 0 0
0
0
9 2-In AND~
219 423 456 0 3 22
0 6 17 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -591757727
65 0 0 0 4 1 8 0
1 U
9914 0 0
0
0
8 2-In OR~
219 704 472 0 3 22
0 16 15 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -759529873
65 0 0 0 4 1 7 0
1 U
3747 0 0
0
0
9 Inverter~
13 870 525 0 2 22
0 6 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U11B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 6 0
1 U
3549 0 0
0
0
9 Inverter~
13 354 464 0 2 22
0 7 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U11A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 6 0
1 U
7931 0 0
0
0
9 2-In XOR~
219 882 375 0 3 22
0 16 9 21
0
0 0 624 692
6 74LS86
-21 -24 21 -16
4 U10A
-10 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
9325 0 0
0
0
9 2-In XOR~
219 883 417 0 3 22
0 18 9 22
0
0 0 624 692
6 74LS86
-21 -24 21 -16
3 U7D
-7 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 4 0
1 U
8903 0 0
0
0
9 2-In XOR~
219 880 333 0 3 22
0 15 9 20
0
0 0 624 692
6 74LS86
-21 -24 21 -16
3 U7C
-7 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 4 0
1 U
3834 0 0
0
0
9 2-In XOR~
219 879 291 0 3 22
0 13 9 19
0
0 0 624 692
6 74LS86
-21 -24 21 -16
3 U7B
-7 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 4 0
1 U
3363 0 0
0
0
7 Ground~
168 987 494 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7668 0 0
0
0
6 74LS47
187 1070 298 0 14 29
0 33 32 31 30 57 58 23 24 25
26 27 28 29 59
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U9
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
6 74LS83
105 1029 415 0 14 29
0 19 20 21 22 2 3 3 2 9
33 32 31 30 60
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3874 0 0
0
0
2 +V
167 981 58 0 1 3
0 34
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6671 0 0
0
0
9 CA 7-Seg~
184 1034 156 0 18 19
10 29 28 27 26 25 24 23 61 34
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3789 0 0
0
0
9 CA 7-Seg~
184 935 157 0 18 19
10 62 4 4 63 64 65 5 66 34
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4871 0 0
0
0
9 2-In XOR~
219 271 282 0 3 22
0 6 38 42
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3750 0 0
0
0
9 2-In XOR~
219 341 281 0 3 22
0 6 35 41
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
8778 0 0
0
0
9 2-In XOR~
219 406 284 0 3 22
0 6 36 40
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
538 0 0
0
0
9 2-In XOR~
219 476 283 0 3 22
0 6 37 39
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
6843 0 0
0
0
6 74LS83
105 525 388 0 14 29
0 43 44 45 46 39 40 41 42 6
13 15 16 18 7
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3136 0 0
0
0
14 Logic Display~
6 633 78 0 1 2
10 43
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5950 0 0
0
0
14 Logic Display~
6 667 77 0 1 2
10 44
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 702 77 0 1 2
10 45
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 734 78 0 1 2
10 46
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
7 Ground~
168 487 227 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
7 74LS173
129 529 145 0 14 29
0 2 2 2 47 48 6 49 50 2
2 43 44 45 46
0
0 0 13040 692
7 74LS173
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4132 0 0
0
0
14 Logic Display~
6 460 34 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4551 0 0
0
0
14 Logic Display~
6 426 35 0 1 2
10 35
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3635 0 0
0
0
14 Logic Display~
6 391 35 0 1 2
10 36
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3973 0 0
0
0
14 Logic Display~
6 357 36 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3851 0 0
0
0
2 +V
167 225 201 0 1 3
0 51
0
0 0 54256 180
2 5V
7 -2 21 6
2 V1
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8383 0 0
0
0
10 Ascii Key~
169 124 97 0 11 12
0 56 55 54 53 67 68 69 52 0
0 55
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
9334 0 0
0
0
7 Buffer~
58 203 149 0 2 22
0 52 47
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
7471 0 0
0
0
7 74LS273
150 263 118 0 18 37
0 51 47 37 36 35 38 53 54 55
56 48 6 49 50 37 36 35 38
0
0 0 13040 692
7 74LS273
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
3334 0 0
0
0
96
1 0 3 0 0 4224 0 1 0 0 15 2
965 280
965 424
3 0 4 0 0 4096 0 20 0 0 3 2
926 193
926 236
2 2 4 0 0 8320 0 20 1 0 0 4
920 193
920 236
965 236
965 244
3 7 5 0 0 4224 0 2 20 0 0 3
840 206
950 206
950 193
1 0 6 0 0 4096 0 2 0 0 7 3
789 197
653 197
653 222
1 0 7 0 0 8192 0 3 0 0 10 3
716 237
663 237
663 499
2 0 6 0 0 8192 0 3 0 0 9 3
716 219
653 219
653 525
2 3 8 0 0 4224 0 2 3 0 0 3
789 215
765 215
765 228
1 0 6 0 0 4224 0 9 0 0 63 3
855 525
285 525
285 351
2 0 7 0 0 4224 0 4 0 0 11 2
828 499
482 499
14 1 7 0 0 0 0 25 10 0 0 4
482 422
482 499
339 499
339 464
9 0 9 0 0 4096 0 17 0 0 28 4
997 460
813 460
813 433
639 433
0 1 2 0 0 4096 0 0 15 44 0 2
987 442
987 488
7 0 3 0 0 0 0 17 0 0 15 2
997 433
947 433
6 3 3 0 0 128 0 17 5 0 0 3
997 424
947 424
947 500
2 2 10 0 0 8320 0 5 9 0 0 4
902 509
897 509
897 525
891 525
3 1 11 0 0 8320 0 4 5 0 0 3
874 490
874 491
902 491
3 1 12 0 0 4224 0 6 4 0 0 2
804 481
828 481
2 0 13 0 0 4096 0 6 0 0 32 3
759 490
586 490
586 422
3 1 14 0 0 4224 0 8 6 0 0 2
737 472
759 472
2 0 15 0 0 4096 0 8 0 0 31 3
691 481
597 481
597 429
1 0 16 0 0 4096 0 8 0 0 30 3
691 463
608 463
608 437
2 2 17 0 0 8320 0 7 10 0 0 3
399 465
399 464
375 464
1 0 6 0 0 0 0 7 0 0 63 2
399 447
399 351
2 0 9 0 0 4224 0 12 0 0 28 2
867 408
639 408
2 0 9 0 0 0 0 11 0 0 28 2
866 366
639 366
2 0 9 0 0 0 0 13 0 0 28 2
864 324
639 324
3 2 9 0 0 0 0 7 14 0 0 5
444 456
444 455
639 455
639 282
863 282
13 1 18 0 0 8320 0 25 12 0 0 4
509 422
509 445
867 445
867 426
12 1 16 0 0 16512 0 25 11 0 0 5
518 422
518 437
628 437
628 384
866 384
11 1 15 0 0 16512 0 25 13 0 0 5
527 422
527 429
620 429
620 342
864 342
10 1 13 0 0 12416 0 25 14 0 0 4
536 422
611 422
611 300
863 300
1 3 19 0 0 8320 0 17 14 0 0 4
997 379
935 379
935 291
912 291
2 3 20 0 0 4224 0 17 13 0 0 4
997 388
926 388
926 333
913 333
3 3 21 0 0 4224 0 17 11 0 0 3
997 397
915 397
915 375
3 4 22 0 0 12416 0 12 17 0 0 4
916 417
932 417
932 406
997 406
7 7 23 0 0 8320 0 16 19 0 0 4
1111 265
1111 216
1049 216
1049 192
6 8 24 0 0 8320 0 19 16 0 0 4
1043 192
1043 223
1102 223
1102 265
9 5 25 0 0 8320 0 16 19 0 0 4
1093 265
1093 228
1037 228
1037 192
4 10 26 0 0 8320 0 19 16 0 0 4
1031 192
1031 233
1084 233
1084 265
11 3 27 0 0 8320 0 16 19 0 0 4
1075 265
1075 239
1025 239
1025 192
2 12 28 0 0 4224 0 19 16 0 0 4
1019 192
1019 243
1066 243
1066 265
13 1 29 0 0 12416 0 16 19 0 0 4
1057 265
1057 248
1013 248
1013 192
5 8 2 0 0 0 0 17 17 0 0 4
997 415
987 415
987 442
997 442
13 4 30 0 0 8320 0 17 16 0 0 3
1061 433
1084 433
1084 335
12 3 31 0 0 8320 0 17 16 0 0 3
1061 424
1093 424
1093 335
11 2 32 0 0 8320 0 17 16 0 0 3
1061 415
1102 415
1102 335
1 10 33 0 0 4224 0 16 17 0 0 3
1111 335
1111 406
1061 406
9 0 34 0 0 8320 0 19 0 0 50 3
1034 120
1034 92
980 92
9 1 34 0 0 0 0 20 18 0 0 4
935 121
935 92
981 92
981 67
2 0 35 0 0 4096 0 22 0 0 84 4
353 262
353 173
335 173
335 86
2 0 36 0 0 4224 0 23 0 0 83 3
418 265
418 95
386 95
2 0 37 0 0 12416 0 24 0 0 82 5
488 264
488 242
445 242
445 103
357 103
2 0 38 0 0 12288 0 21 0 0 85 4
283 263
283 186
323 186
323 77
5 3 39 0 0 8320 0 25 24 0 0 4
527 358
527 322
479 322
479 313
3 6 40 0 0 8320 0 23 25 0 0 4
409 314
409 332
518 332
518 358
7 3 41 0 0 8320 0 25 22 0 0 4
509 358
509 338
344 338
344 311
3 8 42 0 0 8320 0 21 25 0 0 4
274 312
274 345
500 345
500 358
1 0 6 0 0 0 0 21 0 0 62 2
265 263
265 253
1 0 6 0 0 0 0 24 0 0 61 3
470 264
470 253
400 253
1 0 6 0 0 0 0 23 0 0 62 3
400 265
400 253
335 253
1 0 6 0 0 0 0 22 0 0 63 3
335 262
335 253
247 253
9 0 6 0 0 128 0 25 0 0 79 6
482 358
482 351
247 351
247 179
303 179
303 131
1 0 43 0 0 12416 0 25 0 0 68 4
563 358
563 286
623 286
623 140
2 0 44 0 0 12416 0 25 0 0 69 4
554 358
554 279
612 279
612 131
3 0 45 0 0 12416 0 25 0 0 70 4
545 358
545 268
603 268
603 122
4 0 46 0 0 12288 0 25 0 0 71 4
536 358
536 260
593 260
593 113
11 1 43 0 0 0 0 31 26 0 0 3
561 140
633 140
633 96
12 1 44 0 0 0 0 31 27 0 0 3
561 131
667 131
667 95
13 1 45 0 0 0 0 31 28 0 0 3
561 122
702 122
702 95
14 1 46 0 0 4224 0 31 29 0 0 3
561 113
734 113
734 96
2 4 47 0 0 8320 0 38 31 0 0 5
218 149
218 217
479 217
479 149
497 149
2 0 2 0 0 0 0 31 0 0 75 2
491 167
487 167
1 0 2 0 0 0 0 31 0 0 75 2
497 176
487 176
3 0 2 0 0 8192 0 31 0 0 77 3
491 158
487 158
487 205
9 0 2 0 0 0 0 31 0 0 77 2
567 176
580 176
10 1 2 0 0 12416 0 31 30 0 0 5
567 167
580 167
580 205
487 205
487 221
11 5 48 0 0 4224 0 39 31 0 0 2
295 140
497 140
12 6 6 0 0 0 0 39 31 0 0 2
295 131
497 131
13 7 49 0 0 4224 0 39 31 0 0 2
295 122
497 122
14 8 50 0 0 4224 0 39 31 0 0 2
295 113
497 113
1 15 37 0 0 0 0 35 39 0 0 3
357 54
357 104
295 104
1 16 36 0 0 0 0 34 39 0 0 3
391 53
391 95
295 95
1 17 35 0 0 8320 0 33 39 0 0 3
426 53
426 86
295 86
1 18 38 0 0 8320 0 32 39 0 0 3
460 52
460 77
295 77
17 5 35 0 0 0 0 39 39 0 0 6
295 86
303 86
303 31
206 31
206 122
231 122
4 16 36 0 0 0 0 39 39 0 0 6
231 131
219 131
219 20
310 20
310 95
295 95
3 15 37 0 0 0 0 39 39 0 0 6
231 140
223 140
223 15
317 15
317 104
295 104
18 6 38 0 0 0 0 39 39 0 0 5
295 77
295 49
212 49
212 113
231 113
1 1 51 0 0 4224 0 39 36 0 0 2
225 158
225 186
2 2 47 0 0 0 0 38 39 0 0 2
218 149
231 149
8 1 52 0 0 8320 0 37 38 0 0 4
149 117
180 117
180 149
188 149
4 7 53 0 0 4224 0 37 39 0 0 4
149 93
217 93
217 104
231 104
3 8 54 0 0 4224 0 37 39 0 0 4
149 87
217 87
217 95
231 95
2 9 55 0 0 4224 0 37 39 0 0 4
149 81
217 81
217 86
231 86
1 10 56 0 0 4224 0 37 39 0 0 4
149 75
217 75
217 77
231 77
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
