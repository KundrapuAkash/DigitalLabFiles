CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 1061 291 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1063 339 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 711 160 0 1 2
10 5
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 740 160 0 1 2
10 6
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 769 160 0 1 2
10 7
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 798 160 0 1 2
10 8
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 592 410 0 1 2
10 13
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 563 410 0 1 2
10 14
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 534 410 0 1 2
10 15
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 505 410 0 1 2
10 16
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 712 410 0 1 2
10 9
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 683 410 0 1 2
10 10
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 654 410 0 1 2
10 11
0
0 0 53856 512
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 625 410 0 1 2
10 12
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
2 +V
167 937 292 0 1 3
0 17
0
0 0 54256 180
2 5V
7 -2 21 6
2 V2
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
7 Ground~
168 1053 255 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
14 Logic Display~
6 1002 87 0 1 2
10 21
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 973 87 0 1 2
10 20
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 944 87 0 1 2
10 19
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 915 87 0 1 2
10 18
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 450 27 0 1 2
10 25
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 479 27 0 1 2
10 24
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 508 27 0 1 2
10 23
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 537 27 0 1 2
10 22
0
0 0 53856 512
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6843 0 0
0
0
10 Ascii Key~
169 1057 148 0 11 12
0 21 20 19 18 42 43 44 45 0
0 51
0
0 0 4656 602
0
4 KBD2
-12 -39 16 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3136 0 0
0
0
7 74LS193
137 889 233 0 14 29
0 17 4 3 2 18 19 20 21 46
47 5 6 7 8
0
0 0 13040 180
7 74LS193
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
5950 0 0
0
0
2 +V
167 243 330 0 1 3
0 26
0
0 0 54256 90
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5670 0 0
0
0
7 74LS273
150 331 361 0 18 37
0 26 4 27 28 29 30 31 32 33
34 16 15 14 13 12 11 10 9
0
0 0 13040 782
7 74LS273
-24 -60 25 -52
2 U5
54 0 68 8
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
6828 0 0
0
0
7 Ground~
168 432 206 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6735 0 0
0
0
7 Ground~
168 289 204 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8365 0 0
0
0
6 74LS83
105 355 239 0 14 29
0 12 11 10 9 25 24 23 22 2
31 32 33 34 35
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4132 0 0
0
0
6 74LS83
105 225 238 0 14 29
0 16 15 14 13 2 2 2 2 35
27 28 29 30 48
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U2
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4551 0 0
0
0
7 Buffer~
58 114 62 0 2 22
0 41 40
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3635 0 0
0
0
10 Ascii Key~
169 50 42 0 11 12
0 39 38 37 36 49 50 51 41 0
0 53
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3973 0 0
0
0
7 74LS173
129 188 57 0 14 29
0 2 2 2 40 36 37 38 39 2
2 25 24 23 22
0
0 0 13040 692
7 74LS173
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3851 0 0
0
0
7 Ground~
168 137 120 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8383 0 0
0
0
67
3 1 3 0 0 4224 0 26 1 0 0 4
927 246
1020 246
1020 291
1049 291
2 0 4 0 0 8320 0 28 0 0 3 3
299 334
299 318
1010 318
2 1 4 0 0 0 0 26 2 0 0 4
921 255
1010 255
1010 339
1051 339
11 1 5 0 0 4224 0 26 3 0 0 3
857 228
711 228
711 178
12 1 6 0 0 4224 0 26 4 0 0 3
857 219
740 219
740 178
13 1 7 0 0 4224 0 26 5 0 0 3
857 210
769 210
769 178
14 1 8 0 0 4224 0 26 6 0 0 3
857 201
798 201
798 178
0 1 9 0 0 8320 0 0 11 30 0 4
238 476
238 519
712 519
712 428
0 1 10 0 0 8320 0 0 12 31 0 4
244 467
244 514
683 514
683 428
0 1 11 0 0 8320 0 0 13 32 0 4
250 457
250 510
654 510
654 428
0 1 12 0 0 8320 0 0 14 33 0 4
260 445
260 505
625 505
625 428
0 1 13 0 0 8320 0 0 7 34 0 4
268 435
268 500
592 500
592 428
0 1 14 0 0 8320 0 0 8 35 0 4
277 426
277 495
563 495
563 428
0 1 15 0 0 8320 0 0 9 36 0 4
286 417
286 489
534 489
534 428
0 1 16 0 0 8320 0 0 10 37 0 4
295 408
295 483
505 483
505 428
1 1 17 0 0 4224 0 26 15 0 0 3
921 264
937 264
937 277
4 1 2 0 0 4224 0 26 16 0 0 3
921 237
1053 237
1053 249
0 5 18 0 0 4096 0 0 26 22 0 3
933 144
933 228
921 228
0 6 19 0 0 4096 0 0 26 23 0 3
963 138
963 219
921 219
0 7 20 0 0 4224 0 0 26 24 0 3
993 132
993 210
921 210
0 8 21 0 0 8320 0 0 26 25 0 3
1016 126
1016 201
921 201
4 1 18 0 0 4224 0 25 20 0 0 3
1032 144
915 144
915 105
3 1 19 0 0 4224 0 25 19 0 0 3
1032 138
944 138
944 105
2 1 20 0 0 0 0 25 18 0 0 3
1032 132
973 132
973 105
1 1 21 0 0 0 0 25 17 0 0 3
1032 126
1002 126
1002 105
1 0 22 0 0 8192 0 24 0 0 52 3
537 45
537 84
380 84
1 0 23 0 0 8192 0 23 0 0 51 3
508 45
508 73
371 73
1 0 24 0 0 8192 0 22 0 0 50 3
479 45
479 62
362 62
1 0 25 0 0 8192 0 21 0 0 49 3
450 45
450 52
353 52
4 18 9 0 0 0 0 31 28 0 0 6
344 209
344 132
73 132
73 476
371 476
371 398
17 3 10 0 0 0 0 28 31 0 0 6
362 398
362 467
87 467
87 143
335 143
335 209
16 2 11 0 0 0 0 28 31 0 0 6
353 398
353 457
100 457
100 156
326 156
326 209
15 1 12 0 0 0 0 28 31 0 0 6
344 398
344 445
112 445
112 168
317 168
317 209
4 14 13 0 0 0 0 32 28 0 0 6
214 208
214 179
124 179
124 435
335 435
335 398
13 3 14 0 0 0 0 28 32 0 0 6
326 398
326 426
137 426
137 189
205 189
205 208
12 2 15 0 0 0 0 28 32 0 0 6
317 398
317 417
147 417
147 198
196 198
196 208
11 1 16 0 0 0 0 28 32 0 0 5
308 398
308 408
158 408
158 208
187 208
1 1 26 0 0 4224 0 28 27 0 0 2
290 328
254 328
10 3 27 0 0 8320 0 32 28 0 0 4
214 272
214 303
308 303
308 334
11 4 28 0 0 8320 0 32 28 0 0 4
223 272
223 295
317 295
317 334
12 5 29 0 0 8320 0 32 28 0 0 4
232 272
232 287
326 287
326 334
13 6 30 0 0 8320 0 32 28 0 0 4
241 272
241 279
335 279
335 334
10 7 31 0 0 4224 0 31 28 0 0 2
344 273
344 334
11 8 32 0 0 4224 0 31 28 0 0 2
353 273
353 334
12 9 33 0 0 4224 0 31 28 0 0 2
362 273
362 334
13 10 34 0 0 4224 0 31 28 0 0 2
371 273
371 334
14 9 35 0 0 16512 0 31 32 0 0 6
398 273
398 286
445 286
445 178
268 178
268 208
9 1 2 0 0 0 0 31 29 0 0 4
398 209
398 189
432 189
432 200
11 5 25 0 0 8320 0 35 31 0 0 3
220 52
353 52
353 209
12 6 24 0 0 8320 0 35 31 0 0 3
220 43
362 43
362 209
13 7 23 0 0 8320 0 35 31 0 0 3
220 34
371 34
371 209
14 8 22 0 0 8320 0 35 31 0 0 3
220 25
380 25
380 209
8 0 2 0 0 0 0 32 0 0 56 2
250 208
250 189
7 0 2 0 0 0 0 32 0 0 56 2
241 208
241 189
6 0 2 0 0 0 0 32 0 0 56 2
232 208
232 189
5 1 2 0 0 0 0 32 30 0 0 4
223 208
223 189
289 189
289 198
2 0 2 0 0 0 0 35 0 0 58 2
150 79
137 79
3 1 2 0 0 0 0 35 36 0 0 3
150 70
137 70
137 114
9 0 2 0 0 0 0 35 0 0 60 2
226 88
239 88
10 0 2 0 0 0 0 35 0 0 61 4
226 79
239 79
239 108
137 108
1 1 2 0 0 0 0 35 36 0 0 3
156 88
137 88
137 114
4 5 36 0 0 4224 0 34 35 0 0 4
75 38
142 38
142 52
156 52
3 6 37 0 0 4224 0 34 35 0 0 4
75 32
142 32
142 43
156 43
2 7 38 0 0 4224 0 34 35 0 0 4
75 26
142 26
142 34
156 34
1 8 39 0 0 4224 0 34 35 0 0 4
75 20
142 20
142 25
156 25
2 4 40 0 0 12416 0 33 35 0 0 4
129 62
142 62
142 61
156 61
8 1 41 0 0 4224 0 34 33 0 0 2
75 62
99 62
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
