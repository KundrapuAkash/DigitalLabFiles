CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
24
14 Logic Display~
6 737 374 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 855 374 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 820 374 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 786 375 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 887 375 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
9 2-In XOR~
219 271 282 0 3 22
0 16 11 15
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5D
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 341 281 0 3 22
0 16 8 14
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5C
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 406 284 0 3 22
0 16 9 13
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5A
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
9 2-In XOR~
219 476 283 0 3 22
0 16 10 12
0
0 0 624 782
6 74LS86
-21 -24 21 -16
3 U5B
26 -6 47 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3549 0 0
0
0
6 74LS83
105 525 388 0 14 29
0 17 18 19 20 12 13 14 15 16
4 5 6 7 3
0
0 0 13040 270
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
14 Logic Display~
6 633 78 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 667 77 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 702 77 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 734 78 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
7 Ground~
168 487 227 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7668 0 0
0
0
7 74LS173
129 529 145 0 14 29
0 2 2 2 21 22 16 23 24 2
2 17 18 19 20
0
0 0 13040 692
7 74LS173
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
14 Logic Display~
6 460 34 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 426 35 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 391 35 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 357 36 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
2 +V
167 225 201 0 1 3
0 25
0
0 0 54256 180
2 5V
7 -2 21 6
2 V1
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3750 0 0
0
0
10 Ascii Key~
169 124 97 0 11 12
0 30 29 28 27 31 32 33 26 0
1 32
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
8778 0 0
0
0
7 Buffer~
58 203 149 0 2 22
0 26 21
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
538 0 0
0
0
7 74LS273
150 263 118 0 18 37
0 25 21 10 9 8 11 27 28 29
30 22 16 23 24 10 9 8 11
0
0 0 13040 692
7 74LS273
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
51
1 14 3 0 0 8320 0 1 10 0 0 4
737 392
737 459
482 459
482 422
10 1 4 0 0 4224 0 10 4 0 0 3
536 422
786 422
786 393
11 1 5 0 0 8320 0 10 3 0 0 4
527 422
527 433
820 433
820 392
12 1 6 0 0 8320 0 10 2 0 0 4
518 422
518 441
855 441
855 392
13 1 7 0 0 8320 0 10 5 0 0 4
509 422
509 448
887 448
887 393
2 0 8 0 0 4096 0 7 0 0 39 4
353 262
353 173
335 173
335 86
2 0 9 0 0 4224 0 8 0 0 38 3
418 265
418 95
386 95
2 0 10 0 0 12416 0 9 0 0 37 5
488 264
488 242
445 242
445 103
357 103
2 0 11 0 0 12288 0 6 0 0 40 4
283 263
283 186
323 186
323 77
5 3 12 0 0 8320 0 10 9 0 0 4
527 358
527 322
479 322
479 313
3 6 13 0 0 8320 0 8 10 0 0 4
409 314
409 332
518 332
518 358
7 3 14 0 0 8320 0 10 7 0 0 4
509 358
509 338
344 338
344 311
3 8 15 0 0 8320 0 6 10 0 0 4
274 312
274 345
500 345
500 358
1 0 16 0 0 4096 0 6 0 0 17 2
265 263
265 253
1 0 16 0 0 8192 0 9 0 0 16 3
470 264
470 253
400 253
1 0 16 0 0 0 0 8 0 0 17 3
400 265
400 253
335 253
1 0 16 0 0 8192 0 7 0 0 18 3
335 262
335 253
247 253
9 0 16 0 0 8320 0 10 0 0 34 6
482 358
482 351
247 351
247 179
303 179
303 131
1 0 17 0 0 12416 0 10 0 0 23 4
563 358
563 286
623 286
623 140
2 0 18 0 0 12416 0 10 0 0 24 4
554 358
554 279
612 279
612 131
3 0 19 0 0 12416 0 10 0 0 25 4
545 358
545 268
603 268
603 122
4 0 20 0 0 12288 0 10 0 0 26 4
536 358
536 260
593 260
593 113
11 1 17 0 0 128 0 16 11 0 0 3
561 140
633 140
633 96
12 1 18 0 0 128 0 16 12 0 0 3
561 131
667 131
667 95
13 1 19 0 0 128 0 16 13 0 0 3
561 122
702 122
702 95
14 1 20 0 0 4224 0 16 14 0 0 3
561 113
734 113
734 96
2 4 21 0 0 8320 0 23 16 0 0 5
218 149
218 217
479 217
479 149
497 149
2 0 2 0 0 4096 0 16 0 0 30 2
491 167
487 167
1 0 2 0 0 4096 0 16 0 0 30 2
497 176
487 176
3 0 2 0 0 8192 0 16 0 0 32 3
491 158
487 158
487 205
9 0 2 0 0 0 0 16 0 0 32 2
567 176
580 176
10 1 2 0 0 12416 0 16 15 0 0 5
567 167
580 167
580 205
487 205
487 221
11 5 22 0 0 4224 0 24 16 0 0 2
295 140
497 140
12 6 16 0 0 128 0 24 16 0 0 2
295 131
497 131
13 7 23 0 0 4224 0 24 16 0 0 2
295 122
497 122
14 8 24 0 0 4224 0 24 16 0 0 2
295 113
497 113
1 15 10 0 0 0 0 20 24 0 0 3
357 54
357 104
295 104
1 16 9 0 0 0 0 19 24 0 0 3
391 53
391 95
295 95
1 17 8 0 0 8320 0 18 24 0 0 3
426 53
426 86
295 86
1 18 11 0 0 8320 0 17 24 0 0 3
460 52
460 77
295 77
17 5 8 0 0 0 0 24 24 0 0 6
295 86
303 86
303 31
206 31
206 122
231 122
4 16 9 0 0 128 0 24 24 0 0 6
231 131
219 131
219 20
310 20
310 95
295 95
3 15 10 0 0 128 0 24 24 0 0 6
231 140
223 140
223 15
317 15
317 104
295 104
18 6 11 0 0 0 0 24 24 0 0 5
295 77
295 49
212 49
212 113
231 113
1 1 25 0 0 4224 0 24 21 0 0 2
225 158
225 186
2 2 21 0 0 128 0 23 24 0 0 2
218 149
231 149
8 1 26 0 0 8320 0 22 23 0 0 4
149 117
180 117
180 149
188 149
4 7 27 0 0 4224 0 22 24 0 0 4
149 93
217 93
217 104
231 104
3 8 28 0 0 4224 0 22 24 0 0 4
149 87
217 87
217 95
231 95
2 9 29 0 0 4224 0 22 24 0 0 4
149 81
217 81
217 86
231 86
1 10 30 0 0 4224 0 22 24 0 0 4
149 75
217 75
217 77
231 77
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
