CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 1003 517 0 1 11
0 6
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1004 484 0 1 11
0 7
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 1004 445 0 1 11
0 8
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 1002 404 0 1 11
0 9
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 805 412 0 1 11
0 22
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 807 453 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 807 492 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 806 525 0 1 11
0 19
0
0 0 21360 512
2 0V
-7 -16 7 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 618 414 0 1 11
0 35
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V9
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 620 455 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 620 494 0 1 11
0 33
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 619 527 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 428 529 0 1 11
0 45
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 429 496 0 1 11
0 46
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 429 457 0 1 11
0 47
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7668 0 0
0
0
13 Logic Switch~
5 427 416 0 1 11
0 48
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4718 0 0
0
0
7 Ground~
168 318 380 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3874 0 0
0
0
6 74LS47
187 937 295 0 14 29
0 9 8 7 6 58 4 14 13 12
11 10 15 16 59
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6671 0 0
0
0
9 CA 7-Seg~
184 959 199 0 18 19
10 16 15 10 11 12 13 14 60 17
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3789 0 0
0
0
2 +V
167 959 80 0 1 3
0 18
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V16
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4871 0 0
0
0
2 +V
167 762 88 0 1 3
0 31
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V15
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3750 0 0
0
0
9 CA 7-Seg~
184 762 207 0 18 19
10 29 28 23 24 25 26 27 61 30
2 2 0 0 0 0 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8778 0 0
0
0
6 74LS47
187 740 303 0 14 29
0 22 21 20 19 62 5 27 26 25
24 23 28 29 4
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U3
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
538 0 0
0
0
2 +V
167 575 90 0 1 3
0 44
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V10
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6843 0 0
0
0
9 CA 7-Seg~
184 575 209 0 18 19
10 42 41 36 37 38 39 40 63 43
0 2 0 0 2 0 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3136 0 0
0
0
6 74LS47
187 553 305 0 14 29
0 35 34 33 32 64 3 40 39 38
37 36 41 42 5
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U2
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5950 0 0
0
0
6 74LS47
187 362 307 0 14 29
0 48 47 46 45 65 2 53 52 51
50 49 54 55 3
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
9 CA 7-Seg~
184 384 211 0 18 19
10 55 54 49 50 51 52 53 66 56
2 2 2 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
6828 0 0
0
0
2 +V
167 384 92 0 1 3
0 57
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6735 0 0
0
0
9 Resistor~
219 959 123 0 4 5
0 17 18 0 1
0
0 0 880 90
3 150
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 762 131 0 4 5
0 30 31 0 1
0
0 0 880 90
3 150
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 575 133 0 4 5
0 43 44 0 1
0
0 0 880 90
3 150
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 384 135 0 4 5
0 56 57 0 1
0
0 0 880 90
3 150
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
56
14 6 3 0 0 12416 0 27 26 0 0 6
322 280
322 39
457 39
457 353
513 353
513 342
14 6 4 0 0 12416 0 23 18 0 0 6
700 276
700 38
844 38
844 353
897 353
897 332
14 6 5 0 0 12416 0 26 23 0 0 6
513 278
513 38
662 38
662 353
700 353
700 340
6 1 2 0 0 4224 0 27 17 0 0 4
322 344
322 366
318 366
318 374
4 1 6 0 0 4240 0 18 1 0 0 3
951 332
951 517
991 517
3 1 7 0 0 4240 0 18 2 0 0 3
960 332
960 484
992 484
2 1 8 0 0 4240 0 18 3 0 0 3
969 332
969 445
992 445
1 1 9 0 0 4240 0 18 4 0 0 3
978 332
978 404
990 404
3 11 10 0 0 4240 0 19 18 0 0 4
950 235
950 249
942 249
942 262
4 10 11 0 0 4240 0 19 18 0 0 4
956 235
956 254
951 254
951 262
5 9 12 0 0 4240 0 19 18 0 0 4
962 235
962 254
960 254
960 262
6 8 13 0 0 8336 0 19 18 0 0 3
968 235
969 235
969 262
7 7 14 0 0 12432 0 19 18 0 0 4
974 235
974 240
978 240
978 262
2 12 15 0 0 12432 0 19 18 0 0 4
944 235
944 243
933 243
933 262
1 13 16 0 0 8336 0 19 18 0 0 3
938 235
924 235
924 262
1 9 17 0 0 4240 0 30 19 0 0 2
959 141
959 163
1 2 18 0 0 4240 0 20 30 0 0 2
959 89
959 105
4 1 19 0 0 4224 0 23 8 0 0 3
754 340
754 525
794 525
3 1 20 0 0 4224 0 23 7 0 0 3
763 340
763 492
795 492
2 1 21 0 0 4224 0 23 6 0 0 3
772 340
772 453
795 453
1 1 22 0 0 4224 0 23 5 0 0 3
781 340
781 412
793 412
3 11 23 0 0 4224 0 22 23 0 0 4
753 243
753 257
745 257
745 270
4 10 24 0 0 4224 0 22 23 0 0 4
759 243
759 262
754 262
754 270
5 9 25 0 0 4224 0 22 23 0 0 4
765 243
765 262
763 262
763 270
6 8 26 0 0 8320 0 22 23 0 0 3
771 243
772 243
772 270
7 7 27 0 0 12416 0 22 23 0 0 4
777 243
777 248
781 248
781 270
2 12 28 0 0 12416 0 22 23 0 0 4
747 243
747 251
736 251
736 270
1 13 29 0 0 8320 0 22 23 0 0 3
741 243
727 243
727 270
1 9 30 0 0 4224 0 31 22 0 0 2
762 149
762 171
1 2 31 0 0 4224 0 21 31 0 0 2
762 97
762 113
4 1 32 0 0 4224 0 26 12 0 0 3
567 342
567 527
607 527
3 1 33 0 0 4224 0 26 11 0 0 3
576 342
576 494
608 494
2 1 34 0 0 4224 0 26 10 0 0 3
585 342
585 455
608 455
1 1 35 0 0 4224 0 26 9 0 0 3
594 342
594 414
606 414
3 11 36 0 0 4224 0 25 26 0 0 4
566 245
566 259
558 259
558 272
4 10 37 0 0 4224 0 25 26 0 0 4
572 245
572 264
567 264
567 272
5 9 38 0 0 4224 0 25 26 0 0 4
578 245
578 264
576 264
576 272
6 8 39 0 0 8320 0 25 26 0 0 3
584 245
585 245
585 272
7 7 40 0 0 12416 0 25 26 0 0 4
590 245
590 250
594 250
594 272
2 12 41 0 0 12416 0 25 26 0 0 4
560 245
560 253
549 253
549 272
1 13 42 0 0 8320 0 25 26 0 0 3
554 245
540 245
540 272
1 9 43 0 0 4224 0 32 25 0 0 2
575 151
575 173
1 2 44 0 0 4224 0 24 32 0 0 2
575 99
575 115
4 1 45 0 0 4224 0 27 13 0 0 3
376 344
376 529
416 529
3 1 46 0 0 4224 0 27 14 0 0 3
385 344
385 496
417 496
2 1 47 0 0 4224 0 27 15 0 0 3
394 344
394 457
417 457
1 1 48 0 0 4224 0 27 16 0 0 3
403 344
403 416
415 416
3 11 49 0 0 4224 0 28 27 0 0 4
375 247
375 261
367 261
367 274
4 10 50 0 0 4224 0 28 27 0 0 4
381 247
381 266
376 266
376 274
5 9 51 0 0 4224 0 28 27 0 0 4
387 247
387 266
385 266
385 274
6 8 52 0 0 8320 0 28 27 0 0 3
393 247
394 247
394 274
7 7 53 0 0 12416 0 28 27 0 0 4
399 247
399 252
403 252
403 274
2 12 54 0 0 12416 0 28 27 0 0 4
369 247
369 255
358 255
358 274
1 13 55 0 0 8320 0 28 27 0 0 3
363 247
349 247
349 274
1 9 56 0 0 4224 0 33 28 0 0 2
384 153
384 175
1 2 57 0 0 4224 0 29 33 0 0 2
384 101
384 117
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
