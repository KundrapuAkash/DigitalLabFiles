CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 86 325 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 87 263 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
7 Ground~
168 564 345 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 415 509 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 74LS173
129 488 502 0 14 29
0 2 2 2 15 11 14 13 12 2
2 10 9 8 7
0
0 0 13040 782
7 74LS173
-24 -51 25 -43
2 U7
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
5394 0 0
0
0
9 Inverter~
13 215 391 0 2 22
0 17 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
7734 0 0
0
0
14 Logic Display~
6 1016 472 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 931 473 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 961 472 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 989 474 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 898 475 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 813 476 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 843 475 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 871 477 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
6 74LS83
105 492 364 0 14 29
0 10 9 8 7 22 21 20 19 2
14 13 12 16 11
0
0 0 13040 782
7 74LS83A
-24 -60 25 -52
2 U4
57 -2 71 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
14 Logic Display~
6 444 91 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
9 2-In AND~
219 596 194 0 3 22
0 30 3 22
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 1 0
1 U
3874 0 0
0
0
9 2-In AND~
219 656 193 0 3 22
0 29 3 21
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
6671 0 0
0
0
9 2-In AND~
219 713 194 0 3 22
0 28 3 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
3789 0 0
0
0
9 2-In AND~
219 771 194 0 3 22
0 27 3 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
4871 0 0
0
0
6 74LS95
110 387 116 0 12 25
0 18 17 17 26 25 24 23 16 3
4 5 6
0
0 0 13040 0
6 74LS95
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
14 Logic Display~
6 585 37 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 615 36 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 643 38 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 670 36 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3136 0 0
0
0
14 Logic Display~
6 304 48 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5950 0 0
0
0
14 Logic Display~
6 277 50 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 249 48 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 219 49 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
10 Ascii Key~
169 819 126 0 11 12
0 27 28 29 30 31 32 33 34 0
0 111
0
0 0 4656 602
0
4 KBD2
-12 -39 16 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
8365 0 0
0
0
10 Ascii Key~
169 118 169 0 11 12
0 26 25 24 23 35 36 37 38 0
0 111
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
4132 0 0
0
0
53
1 0 2 0 0 4096 0 5 0 0 23 2
459 472
459 457
0 1 3 0 0 8320 0 0 7 44 0 6
455 125
455 243
1092 243
1092 582
1016 582
1016 490
10 1 4 0 0 12416 0 21 10 0 0 7
419 134
441 134
441 255
1080 255
1080 571
989 571
989 492
11 1 5 0 0 12416 0 21 9 0 0 7
419 143
429 143
429 267
1067 267
1067 559
961 559
961 490
12 1 6 0 0 8320 0 21 8 0 0 6
419 152
419 277
1055 277
1055 546
931 546
931 491
1 0 7 0 0 8320 0 11 0 0 19 3
898 493
898 583
522 583
1 0 8 0 0 8320 0 14 0 0 18 3
871 495
871 571
513 571
1 0 9 0 0 8320 0 13 0 0 17 3
843 493
843 559
504 559
1 0 10 0 0 8320 0 12 0 0 16 3
813 494
813 546
495 546
14 5 11 0 0 4224 0 15 5 0 0 4
535 398
535 459
495 459
495 472
12 8 12 0 0 12416 0 15 5 0 0 4
499 398
499 431
522 431
522 472
11 7 13 0 0 4224 0 15 5 0 0 4
490 398
490 437
513 437
513 472
10 6 14 0 0 4224 0 15 5 0 0 4
481 398
481 443
504 443
504 472
2 4 15 0 0 12416 0 6 5 0 0 5
236 391
254 391
254 451
486 451
486 472
13 8 16 0 0 12416 0 15 21 0 0 5
508 398
508 407
336 407
336 152
355 152
1 11 10 0 0 0 0 15 5 0 0 6
454 334
454 323
376 323
376 575
495 575
495 536
12 2 9 0 0 0 0 5 15 0 0 6
504 536
504 588
366 588
366 313
463 313
463 334
13 3 8 0 0 0 0 5 15 0 0 6
513 536
513 597
353 597
353 299
472 299
472 334
14 4 7 0 0 0 0 5 15 0 0 6
522 536
522 607
343 607
343 288
481 288
481 334
9 0 2 0 0 0 0 5 0 0 21 2
459 542
459 549
10 0 2 0 0 12416 0 5 0 0 23 5
468 542
468 549
432 549
432 485
415 485
2 0 2 0 0 0 0 5 0 0 23 2
468 466
468 457
3 1 2 0 0 0 0 5 4 0 0 4
477 466
477 457
415 457
415 503
1 9 2 0 0 0 0 3 15 0 0 4
564 339
564 325
535 325
535 334
1 0 17 0 0 8192 0 6 0 0 27 3
200 391
174 391
174 325
3 0 17 0 0 0 0 21 0 0 27 2
349 107
327 107
1 2 17 0 0 4224 0 1 21 0 0 4
98 325
327 325
327 98
349 98
1 1 18 0 0 4224 0 21 2 0 0 4
355 89
164 89
164 263
99 263
3 8 19 0 0 8320 0 20 15 0 0 4
769 217
769 235
517 235
517 334
3 7 20 0 0 8320 0 19 15 0 0 4
711 217
711 229
508 229
508 334
3 6 21 0 0 8320 0 18 15 0 0 4
654 216
654 223
499 223
499 334
3 5 22 0 0 8320 0 17 15 0 0 3
594 217
490 217
490 334
7 0 23 0 0 4224 0 21 0 0 40 2
355 143
219 143
6 0 24 0 0 4224 0 21 0 0 39 2
355 134
249 134
5 0 25 0 0 4096 0 21 0 0 36 2
355 125
277 125
1 2 25 0 0 8320 0 27 31 0 0 3
277 68
277 153
143 153
4 0 26 0 0 8192 0 21 0 0 38 3
355 116
355 117
304 117
1 1 26 0 0 4224 0 31 26 0 0 3
143 147
304 147
304 66
3 1 24 0 0 0 0 31 28 0 0 3
143 159
249 159
249 66
4 1 23 0 0 0 0 31 29 0 0 3
143 165
219 165
219 67
2 0 3 0 0 0 0 17 0 0 44 2
585 172
585 151
2 0 3 0 0 0 0 18 0 0 44 2
645 171
645 151
2 0 3 0 0 0 0 19 0 0 44 2
702 172
702 151
9 2 3 0 0 128 0 21 20 0 0 5
419 125
561 125
561 151
760 151
760 172
1 0 27 0 0 4096 0 20 0 0 53 2
778 172
778 104
1 0 28 0 0 4096 0 19 0 0 52 2
720 172
720 110
1 0 29 0 0 4096 0 18 0 0 51 2
663 171
663 116
1 0 30 0 0 4096 0 17 0 0 50 2
603 172
603 122
1 9 3 0 0 0 0 16 21 0 0 3
444 109
444 125
419 125
4 1 30 0 0 4224 0 30 22 0 0 3
794 122
585 122
585 55
3 1 29 0 0 4224 0 30 23 0 0 3
794 116
615 116
615 54
2 1 28 0 0 4224 0 30 24 0 0 3
794 110
643 110
643 56
1 1 27 0 0 8320 0 25 30 0 0 3
670 54
670 104
794 104
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
