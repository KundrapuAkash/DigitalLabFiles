CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 4 100 9
5 81 1527 809
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
5 81 1527 809
143654930 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 341 366 0 1 11
0 25
0
0 0 21360 0
2 0V
-8 -15 6 -7
2 V6
-9 -25 5 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 290 475 0 1 11
0 28
0
0 0 21360 0
2 0V
-8 -15 6 -7
2 V3
-9 -25 5 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 187 468 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 756 286 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 512
2 5V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
7 Ground~
168 479 373 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
10 2-In NAND~
219 557 209 0 3 22
0 5 4 6
0
0 0 624 90
6 74LS00
-14 -24 28 -16
3 U8A
19 -2 40 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7734 0 0
0
0
2 +V
167 573 56 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
9 CA 7-Seg~
184 662 118 0 18 19
10 6 12 11 10 9 8 7 31 3
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3747 0 0
0
0
6 1K RAM
79 560 367 0 20 41
0 2 2 2 2 2 2 2 24 23
22 32 33 34 35 4 5 14 13 2
15
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
6 74LS93
109 433 403 0 8 17
0 25 25 36 26 24 23 22 37
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
7 Pulser~
4 186 398 0 10 12
0 38 39 30 40 0 0 5 5 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9325 0 0
0
0
9 2-In AND~
219 282 398 0 3 22
0 30 29 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8903 0 0
0
0
8 2-In OR~
219 343 421 0 3 22
0 27 28 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3834 0 0
0
0
7 Ground~
168 906 314 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
7 Buffer~
58 896 367 0 2 22
0 16 21
0
0 0 624 180
4 4050
-14 -19 14 -11
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 3 0
1 U
7668 0 0
0
0
7 74LS173
129 770 376 0 14 29
0 2 2 2 21 17 18 19 20 15
15 4 5 14 13
0
0 0 13040 512
7 74LS173
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
10 Ascii Key~
169 1017 389 0 11 12
0 20 19 18 17 41 42 43 16 0
1 51
0
0 0 4656 270
0
4 KBD1
-12 -38 16 -30
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3874 0 0
0
0
6 74LS47
187 675 256 0 14 29
0 4 5 14 13 44 45 7 8 9
10 11 12 6 46
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
2 U7
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6671 0 0
0
0
49
9 1 3 0 0 8320 0 8 7 0 0 3
662 82
662 65
573 65
19 0 2 0 0 8320 0 9 0 0 9 4
598 331
598 288
490 288
490 321
1 0 2 0 0 0 0 9 0 0 9 2
528 331
506 331
2 0 2 0 0 0 0 9 0 0 9 2
528 340
506 340
3 0 2 0 0 0 0 9 0 0 9 2
528 349
506 349
4 0 2 0 0 0 0 9 0 0 9 2
528 358
506 358
5 0 2 0 0 0 0 9 0 0 9 2
528 367
506 367
6 0 2 0 0 0 0 9 0 0 9 2
528 376
506 376
7 1 2 0 0 0 0 9 5 0 0 5
528 385
506 385
506 321
479 321
479 367
2 0 4 0 0 8192 0 6 0 0 23 5
568 233
568 270
610 270
610 300
639 300
1 0 5 0 0 8192 0 6 0 0 22 5
550 233
550 281
602 281
602 306
648 306
3 0 6 0 0 8320 0 6 0 0 19 3
559 182
559 173
641 173
7 7 7 0 0 4224 0 8 18 0 0 4
677 154
677 214
640 214
640 223
6 8 8 0 0 4224 0 8 18 0 0 4
671 154
671 214
649 214
649 223
5 9 9 0 0 4224 0 8 18 0 0 4
665 154
665 214
658 214
658 223
4 10 10 0 0 4224 0 8 18 0 0 4
659 154
659 214
667 214
667 223
3 11 11 0 0 4224 0 8 18 0 0 4
653 154
653 214
676 214
676 223
2 12 12 0 0 4224 0 8 18 0 0 4
647 154
647 214
685 214
685 223
1 13 6 0 0 0 0 8 18 0 0 4
641 154
641 214
694 214
694 223
4 0 13 0 0 4096 0 18 0 0 27 4
667 293
667 397
666 397
666 412
3 0 14 0 0 4096 0 18 0 0 28 4
658 293
658 388
657 388
657 403
2 0 5 0 0 12288 0 18 0 0 29 4
649 293
649 306
648 306
648 394
1 0 4 0 0 12288 0 18 0 0 30 4
640 293
640 300
639 300
639 385
0 20 15 0 0 4224 0 0 9 25 0 4
732 348
606 348
606 340
598 340
0 10 15 0 0 0 0 0 16 26 0 2
732 348
732 358
1 9 15 0 0 0 0 4 16 0 0 3
744 286
732 286
732 349
18 14 13 0 0 4224 0 9 16 0 0 2
592 412
738 412
17 13 14 0 0 4224 0 9 16 0 0 2
592 403
738 403
16 12 5 0 0 4224 0 9 16 0 0 2
592 394
738 394
15 11 4 0 0 4224 0 9 16 0 0 2
592 385
738 385
3 1 2 0 0 0 0 16 14 0 0 5
808 367
819 367
819 301
906 301
906 308
2 1 2 0 0 0 0 16 14 0 0 5
808 358
819 358
819 301
906 301
906 308
1 1 2 0 0 0 0 16 14 0 0 5
802 349
819 349
819 301
906 301
906 308
1 8 16 0 0 8320 0 15 17 0 0 3
911 367
911 368
993 368
4 5 17 0 0 4224 0 17 16 0 0 4
993 392
824 392
824 385
802 385
3 6 18 0 0 4224 0 17 16 0 0 4
993 398
824 398
824 394
802 394
2 7 19 0 0 12416 0 17 16 0 0 4
993 404
978 404
978 403
802 403
1 8 20 0 0 4224 0 17 16 0 0 4
993 410
824 410
824 412
802 412
4 2 21 0 0 12416 0 16 15 0 0 4
802 376
824 376
824 367
881 367
7 10 22 0 0 4224 0 10 9 0 0 2
465 412
528 412
6 9 23 0 0 4224 0 10 9 0 0 2
465 403
528 403
5 8 24 0 0 4224 0 10 9 0 0 2
465 394
528 394
0 2 25 0 0 8192 0 0 10 44 0 3
387 394
387 403
401 403
1 1 25 0 0 12416 0 1 10 0 0 6
353 366
354 366
354 361
387 361
387 394
401 394
3 4 26 0 0 4224 0 13 10 0 0 2
376 421
395 421
3 1 27 0 0 4224 0 12 13 0 0 4
303 398
322 398
322 412
330 412
1 2 28 0 0 12416 0 2 13 0 0 5
302 475
302 474
322 474
322 430
330 430
1 2 29 0 0 8320 0 3 12 0 0 4
199 468
250 468
250 407
258 407
3 1 30 0 0 4224 0 11 12 0 0 2
210 389
258 389
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
