CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 371 355 0 1 11
0 11
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 371 308 0 1 11
0 9
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 370 256 0 1 11
0 12
0
0 0 21360 512
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 1178 305 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
2 +V
167 923 390 0 1 3
0 8
0
0 0 54256 180
2 5V
7 -2 21 6
2 V5
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
9 Inverter~
13 650 319 0 2 22
0 9 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
7734 0 0
0
0
9 2-In AND~
219 633 449 0 3 22
0 17 18 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 2 0
1 U
9914 0 0
0
0
8 2-In OR~
219 624 503 0 3 22
0 17 18 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
3747 0 0
0
0
8 2-In OR~
219 832 475 0 3 22
0 15 16 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
3549 0 0
0
0
9 2-In AND~
219 751 556 0 3 22
0 14 6 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
7931 0 0
0
0
9 2-In XOR~
219 809 241 0 3 22
0 19 6 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
9325 0 0
0
0
9 2-In XOR~
219 726 192 0 3 22
0 17 18 19
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -369718155
65 0 0 0 4 1 1 0
1 U
8903 0 0
0
0
6 74LS74
17 1032 374 0 12 25
0 10 13 8 8 26 27 28 29 6
30 31 32
0
0 0 13040 0
6 74LS74
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
14 Logic Display~
6 237 420 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 262 421 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 291 418 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 316 419 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
2 +V
167 239 615 0 1 3
0 3
0
0 0 54256 180
2 5V
7 -2 21 6
2 V8
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6671 0 0
0
0
7 Ground~
168 240 640 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3789 0 0
0
0
6 74LS95
110 306 533 0 12 25
0 12 9 11 3 2 3 3 7 18
20 21 22
0
0 0 13040 602
6 74LS95
-21 -51 21 -43
2 U2
45 -6 59 2
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
4871 0 0
0
0
2 +V
167 240 228 0 1 3
0 4
0
0 0 54256 180
2 5V
7 -2 21 6
2 V4
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3750 0 0
0
0
7 Ground~
168 244 254 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8778 0 0
0
0
6 74LS95
110 310 147 0 12 25
0 12 9 11 4 2 2 4 5 17
23 24 25
0
0 0 13040 602
6 74LS95
-21 -51 21 -43
2 U1
45 -6 59 2
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
538 0 0
0
0
14 Logic Display~
6 246 37 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 271 38 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
14 Logic Display~
6 325 36 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5950 0 0
0
0
14 Logic Display~
6 300 35 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5670 0 0
0
0
42
4 1 3 0 0 8320 0 20 18 0 0 4
305 564
305 594
239 594
239 600
7 1 4 0 0 8192 0 23 21 0 0 4
282 178
282 207
240 207
240 213
5 1 2 0 0 4096 0 23 22 0 0 4
300 178
300 240
244 240
244 248
6 1 2 0 0 0 0 23 22 0 0 4
291 178
291 240
244 240
244 248
5 1 2 0 0 4224 0 20 19 0 0 4
296 564
296 628
240 628
240 634
7 1 3 0 0 0 0 20 18 0 0 4
278 564
278 594
239 594
239 600
4 1 4 0 0 8320 0 23 21 0 0 4
309 178
309 207
240 207
240 213
6 1 3 0 0 128 0 20 18 0 0 4
287 564
287 594
239 594
239 600
8 3 5 0 0 12416 0 23 11 0 0 7
273 178
225 178
225 7
829 7
829 207
842 207
842 241
2 0 6 0 0 8192 0 11 0 0 21 3
793 250
789 250
789 318
8 0 7 0 0 8320 0 20 0 0 0 6
269 564
269 576
870 576
870 246
845 246
845 241
1 9 6 0 0 8192 0 4 13 0 0 3
1178 323
1178 347
1064 347
4 0 8 0 0 4224 0 13 0 0 14 2
994 365
923 365
3 1 8 0 0 0 0 13 5 0 0 3
994 356
923 356
923 375
1 0 9 0 0 4096 0 6 0 0 41 4
635 319
332 319
332 265
327 265
2 1 10 0 0 8320 0 6 13 0 0 3
671 319
671 338
1000 338
3 0 11 0 0 12416 0 20 0 0 40 5
314 570
314 674
187 674
187 314
318 314
0 2 9 0 0 8320 0 0 20 41 0 5
327 276
176 276
176 699
323 699
323 570
1 0 12 0 0 12416 0 20 0 0 42 5
332 564
332 649
469 649
469 219
336 219
3 2 13 0 0 8320 0 9 13 0 0 4
865 475
986 475
986 347
1000 347
2 9 6 0 0 12416 0 10 13 0 0 6
727 565
723 565
723 318
1078 318
1078 347
1064 347
3 1 14 0 0 4224 0 8 10 0 0 4
657 503
719 503
719 547
727 547
3 1 15 0 0 4224 0 7 9 0 0 4
654 449
811 449
811 466
819 466
3 2 16 0 0 8320 0 10 9 0 0 4
772 556
811 556
811 484
819 484
1 0 17 0 0 8192 0 8 0 0 31 3
611 494
551 494
551 183
2 0 18 0 0 4096 0 8 0 0 30 3
611 512
350 512
350 457
2 0 18 0 0 0 0 7 0 0 30 4
609 458
409 458
409 454
404 454
1 0 17 0 0 0 0 7 0 0 31 3
609 440
535 440
535 183
3 1 19 0 0 8320 0 12 11 0 0 4
759 192
785 192
785 232
793 232
2 0 18 0 0 4224 0 12 0 0 32 4
710 201
404 201
404 457
316 457
1 0 17 0 0 4224 0 12 0 0 36 4
710 183
355 183
355 84
325 84
1 9 18 0 0 0 0 17 20 0 0 4
316 437
316 492
296 492
296 500
1 10 20 0 0 4224 0 16 20 0 0 4
291 436
291 492
287 492
287 500
1 11 21 0 0 4224 0 15 20 0 0 4
262 439
262 492
278 492
278 500
1 12 22 0 0 4224 0 14 20 0 0 4
237 438
237 492
269 492
269 500
1 9 17 0 0 0 0 26 23 0 0 4
325 54
325 106
300 106
300 114
1 10 23 0 0 4224 0 27 23 0 0 4
300 53
300 106
291 106
291 114
1 11 24 0 0 4224 0 25 23 0 0 4
271 56
271 106
282 106
282 114
1 12 25 0 0 4224 0 24 23 0 0 4
246 55
246 106
273 106
273 114
3 1 11 0 0 0 0 23 1 0 0 3
318 184
318 355
359 355
2 1 9 0 0 0 0 23 2 0 0 3
327 184
327 308
359 308
1 1 12 0 0 0 0 23 3 0 0 3
336 178
336 256
358 256
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
