CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
16
9 Inverter~
13 503 545 0 2 22
0 4 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 4 0
1 U
8953 0 0
0
0
9 Inverter~
13 503 479 0 2 22
0 3 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
4441 0 0
0
0
10 3-In NAND~
219 748 515 0 4 22
0 6 7 5 8
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
3618 0 0
0
0
10 2-In NAND~
219 557 416 0 3 22
0 11 9 10
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6153 0 0
0
0
10 2-In NAND~
219 556 134 0 3 22
0 12 13 18
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
5394 0 0
0
0
10 2-In NAND~
219 557 229 0 3 22
0 13 15 17
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 2088094389
65 0 0 0 4 1 2 0
1 U
7734 0 0
0
0
10 4-In NAND~
219 562 323 0 5 22
0 11 12 13 14 16
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 2088094389
65 0 0 0 2 1 1 0
1 U
9914 0 0
0
0
2 +V
167 213 182 0 1 3
0 19
0
0 0 54256 90
2 5V
-7 -15 7 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3747 0 0
0
0
7 Ground~
168 264 212 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
7 74LS138
19 316 141 0 14 29
0 4 7 3 19 2 2 11 15 28
9 12 13 29 14
0
0 0 13296 0
7 74LS138
-25 -61 24 -53
2 U3
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
2 +V
167 923 58 0 1 3
0 26
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
9 CA 7-Seg~
184 923 133 0 18 19
10 8 20 21 22 23 24 25 30 26
0 0 2 0 0 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8903 0 0
0
0
6 74LS47
187 774 314 0 14 29
0 18 17 16 10 31 32 25 24 23
22 21 20 8 33
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
7 Ground~
168 165 89 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
6 74LS93
109 232 123 0 8 17
0 2 2 34 27 4 7 3 35
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
7 Pulser~
4 129 150 0 10 12
0 36 37 27 38 0 0 5 5 4
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4718 0 0
0
0
37
1 0 3 0 0 8320 0 2 0 0 25 5
488 479
52 479
52 5
279 5
279 132
1 5 4 0 0 8320 0 1 15 0 0 5
488 545
74 545
74 32
264 32
264 114
2 3 5 0 0 4224 0 1 3 0 0 4
524 545
716 545
716 524
724 524
2 1 6 0 0 4224 0 2 3 0 0 4
524 479
716 479
716 506
724 506
0 2 7 0 0 16512 0 0 3 26 0 5
274 123
274 21
64 21
64 515
724 515
4 0 8 0 0 8320 0 3 0 0 7 3
775 515
876 515
876 332
1 13 8 0 0 0 0 12 13 0 0 3
902 169
902 332
812 332
10 2 9 0 0 8320 0 10 4 0 0 4
354 141
481 141
481 425
533 425
3 4 10 0 0 4224 0 4 13 0 0 4
584 416
734 416
734 305
742 305
1 0 11 0 0 4096 0 7 0 0 11 2
538 310
392 310
7 1 11 0 0 8320 0 10 4 0 0 4
354 114
392 114
392 407
533 407
2 0 12 0 0 8320 0 7 0 0 20 3
538 319
432 319
432 150
0 3 13 0 0 4096 0 0 7 21 0 3
424 159
424 328
538 328
14 4 14 0 0 8320 0 10 7 0 0 4
354 177
416 177
416 337
538 337
0 1 13 0 0 0 0 0 6 21 0 3
504 159
504 220
533 220
8 2 15 0 0 4224 0 10 6 0 0 4
354 123
492 123
492 238
533 238
5 3 16 0 0 4224 0 7 13 0 0 4
589 323
722 323
722 296
742 296
3 2 17 0 0 4224 0 6 13 0 0 4
584 229
722 229
722 287
742 287
3 1 18 0 0 4224 0 5 13 0 0 4
583 134
734 134
734 278
742 278
11 1 12 0 0 0 0 10 5 0 0 4
354 150
515 150
515 125
532 125
12 2 13 0 0 4224 0 10 5 0 0 4
354 159
524 159
524 143
532 143
4 1 19 0 0 12416 0 10 8 0 0 4
284 159
256 159
256 180
224 180
6 0 2 0 0 4096 0 10 0 0 24 2
278 177
264 177
1 5 2 0 0 4096 0 9 10 0 0 3
264 206
264 168
278 168
7 3 3 0 0 128 0 15 10 0 0 2
264 132
284 132
6 2 7 0 0 128 0 15 10 0 0 2
264 123
284 123
5 1 4 0 0 128 0 15 10 0 0 2
264 114
284 114
12 2 20 0 0 8320 0 13 12 0 0 3
812 323
908 323
908 169
11 3 21 0 0 8320 0 13 12 0 0 3
812 314
914 314
914 169
10 4 22 0 0 8320 0 13 12 0 0 3
812 305
920 305
920 169
9 5 23 0 0 8320 0 13 12 0 0 3
812 296
926 296
926 169
8 6 24 0 0 4224 0 13 12 0 0 3
812 287
932 287
932 169
7 7 25 0 0 4224 0 13 12 0 0 3
812 278
938 278
938 169
1 9 26 0 0 4224 0 11 12 0 0 2
923 67
923 97
1 0 2 0 0 4224 0 15 0 0 36 2
200 114
151 114
2 1 2 0 0 0 0 15 14 0 0 5
200 123
151 123
151 75
165 75
165 83
4 3 27 0 0 4224 0 15 16 0 0 2
194 141
153 141
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
