CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 28 100 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 96 1498 799
143654930 0
0
6 Title:
5 Name:
0
0
0
25
7 Ground~
168 784 454 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 575 473 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 405 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 991 472 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
2 +V
167 368 43 0 1 3
0 21
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
6 74LS90
107 385 392 0 10 21
0 2 56 4 3 6 10 11 12 4
10
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U8
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
6 74LS47
187 351 266 0 14 29
0 11 12 4 10 57 58 13 14 15
16 17 18 19 59
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U7
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
9 CA 7-Seg~
184 370 160 0 18 19
10 19 18 17 16 15 14 13 60 20
0 0 0 0 0 0 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3747 0 0
0
0
9 CA 7-Seg~
184 550 164 0 18 19
10 30 29 28 27 26 25 24 61 31
0 0 0 0 2 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
6 74LS47
187 531 270 0 14 29
0 6 3 23 22 62 63 24 25 26
27 28 29 30 64
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U6
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
6 74LS90
107 565 396 0 10 21
0 2 65 4 3 5 22 6 3 23
22
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U5
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
2 +V
167 548 47 0 1 3
0 32
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8903 0 0
0
0
2 +V
167 747 52 0 1 3
0 43
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3834 0 0
0
0
6 74LS90
107 764 401 0 10 21
0 2 66 5 7 8 33 34 5 7
33
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U4
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
6 74LS47
187 730 275 0 14 29
0 34 5 7 33 67 68 35 36 37
38 39 40 41 69
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U3
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
9 CA 7-Seg~
184 749 169 0 18 19
10 41 40 39 38 37 36 35 70 42
0 0 2 0 0 2 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4718 0 0
0
0
9 CA 7-Seg~
184 964 170 0 18 19
10 53 52 51 50 49 48 47 71 54
0 0 0 2 2 2 2 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3874 0 0
0
0
6 74LS47
187 945 276 0 14 29
0 8 45 46 44 72 73 47 48 49
50 51 52 53 74
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6671 0 0
0
0
6 74LS90
107 979 402 0 10 21
0 2 75 2 76 9 44 8 45 46
44
0
0 0 13040 602
6 74LS90
-21 -51 21 -43
2 U2
40 -11 54 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
0
0
2 +V
167 962 53 0 1 3
0 55
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4871 0 0
0
0
7 Pulser~
4 914 537 0 10 12
0 77 78 9 79 0 0 5 5 2
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3750 0 0
0
0
9 Resistor~
219 367 81 0 3 5
0 21 20 1
0
0 0 880 782
3 150
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 547 85 0 3 5
0 32 31 1
0
0 0 880 782
3 150
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 746 90 0 3 5
0 43 42 1
0
0 0 880 782
3 150
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 961 91 0 3 5
0 55 54 1
0
0 0 880 782
3 150
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
71
4 0 3 0 0 8192 0 6 0 0 3 5
379 418
379 469
491 469
491 381
500 381
3 0 4 0 0 8192 0 11 0 0 10 3
568 422
568 455
445 455
4 0 3 0 0 12416 0 11 0 0 32 5
559 422
559 448
500 448
500 333
560 333
5 0 5 0 0 8320 0 11 0 0 46 5
541 428
541 531
824 531
824 340
759 340
3 0 5 0 0 128 0 14 0 0 46 5
767 427
767 471
687 471
687 328
759 328
1 1 2 0 0 4096 0 14 1 0 0 4
785 427
785 440
784 440
784 448
1 1 2 0 0 4224 0 11 2 0 0 4
586 422
586 459
575 459
575 467
5 0 6 0 0 8320 0 6 0 0 31 5
361 424
361 603
628 603
628 336
586 336
1 1 2 0 0 0 0 6 3 0 0 4
406 418
406 429
405 429
405 435
3 0 4 0 0 12416 0 6 0 0 19 5
388 418
388 455
450 455
450 324
370 324
4 0 7 0 0 12416 0 14 0 0 47 5
758 427
758 466
699 466
699 337
749 337
5 7 8 0 0 8320 0 14 19 0 0 5
740 433
740 604
1042 604
1042 364
1000 364
3 0 2 0 0 0 0 19 0 0 14 4
982 428
982 453
994 453
994 458
1 1 2 0 0 0 0 19 4 0 0 4
1000 428
1000 458
991 458
991 466
3 5 9 0 0 8320 0 21 19 0 0 3
938 528
955 528
955 434
10 6 10 0 0 12416 0 6 6 0 0 6
352 354
352 350
338 350
338 432
352 432
352 424
1 7 11 0 0 8320 0 7 6 0 0 3
392 303
406 303
406 354
2 8 12 0 0 8320 0 7 6 0 0 5
383 303
380 303
380 346
388 346
388 354
3 9 4 0 0 0 0 7 6 0 0 3
374 303
370 303
370 354
4 10 10 0 0 0 0 7 6 0 0 3
365 303
352 303
352 354
7 7 13 0 0 12416 0 8 7 0 0 4
385 196
385 207
392 207
392 233
6 8 14 0 0 12416 0 8 7 0 0 4
379 196
379 211
383 211
383 233
5 9 15 0 0 4224 0 8 7 0 0 4
373 196
373 225
374 225
374 233
4 10 16 0 0 4224 0 8 7 0 0 4
367 196
367 225
365 225
365 233
3 11 17 0 0 12416 0 8 7 0 0 4
361 196
361 210
356 210
356 233
2 12 18 0 0 12416 0 8 7 0 0 4
355 196
355 205
347 205
347 233
1 13 19 0 0 8320 0 8 7 0 0 3
349 196
338 196
338 233
2 9 20 0 0 4224 0 22 8 0 0 4
367 99
367 116
370 116
370 124
1 1 21 0 0 12416 0 5 22 0 0 4
368 52
368 57
367 57
367 63
10 6 22 0 0 12416 0 11 11 0 0 6
532 358
532 354
518 354
518 436
532 436
532 428
1 7 6 0 0 0 0 10 11 0 0 3
572 307
586 307
586 358
2 8 3 0 0 128 0 10 11 0 0 5
563 307
560 307
560 350
568 350
568 358
3 9 23 0 0 8320 0 10 11 0 0 3
554 307
550 307
550 358
4 10 22 0 0 0 0 10 11 0 0 3
545 307
532 307
532 358
7 7 24 0 0 12416 0 9 10 0 0 4
565 200
565 211
572 211
572 237
6 8 25 0 0 12416 0 9 10 0 0 4
559 200
559 215
563 215
563 237
5 9 26 0 0 4224 0 9 10 0 0 4
553 200
553 229
554 229
554 237
4 10 27 0 0 4224 0 9 10 0 0 4
547 200
547 229
545 229
545 237
3 11 28 0 0 12416 0 9 10 0 0 4
541 200
541 214
536 214
536 237
2 12 29 0 0 12416 0 9 10 0 0 4
535 200
535 209
527 209
527 237
1 13 30 0 0 8320 0 9 10 0 0 3
529 200
518 200
518 237
2 9 31 0 0 4224 0 23 9 0 0 4
547 103
547 120
550 120
550 128
1 1 32 0 0 12416 0 12 23 0 0 4
548 56
548 61
547 61
547 67
10 6 33 0 0 12416 0 14 14 0 0 6
731 363
731 359
717 359
717 441
731 441
731 433
1 7 34 0 0 8320 0 15 14 0 0 3
771 312
785 312
785 363
2 8 5 0 0 0 0 15 14 0 0 5
762 312
759 312
759 355
767 355
767 363
3 9 7 0 0 0 0 15 14 0 0 3
753 312
749 312
749 363
4 10 33 0 0 0 0 15 14 0 0 3
744 312
731 312
731 363
7 7 35 0 0 12416 0 16 15 0 0 4
764 205
764 216
771 216
771 242
6 8 36 0 0 12416 0 16 15 0 0 4
758 205
758 220
762 220
762 242
5 9 37 0 0 4224 0 16 15 0 0 4
752 205
752 234
753 234
753 242
4 10 38 0 0 4224 0 16 15 0 0 4
746 205
746 234
744 234
744 242
3 11 39 0 0 12416 0 16 15 0 0 4
740 205
740 219
735 219
735 242
2 12 40 0 0 12416 0 16 15 0 0 4
734 205
734 214
726 214
726 242
1 13 41 0 0 8320 0 16 15 0 0 3
728 205
717 205
717 242
2 9 42 0 0 4224 0 24 16 0 0 4
746 108
746 125
749 125
749 133
1 1 43 0 0 12416 0 13 24 0 0 4
747 61
747 66
746 66
746 72
10 6 44 0 0 12416 0 19 19 0 0 6
946 364
946 360
932 360
932 442
946 442
946 434
1 7 8 0 0 0 0 18 19 0 0 3
986 313
1000 313
1000 364
2 8 45 0 0 8320 0 18 19 0 0 5
977 313
974 313
974 356
982 356
982 364
3 9 46 0 0 8320 0 18 19 0 0 3
968 313
964 313
964 364
4 10 44 0 0 0 0 18 19 0 0 3
959 313
946 313
946 364
7 7 47 0 0 12416 0 17 18 0 0 4
979 206
979 217
986 217
986 243
6 8 48 0 0 12416 0 17 18 0 0 4
973 206
973 221
977 221
977 243
5 9 49 0 0 4224 0 17 18 0 0 4
967 206
967 235
968 235
968 243
4 10 50 0 0 4224 0 17 18 0 0 4
961 206
961 235
959 235
959 243
3 11 51 0 0 12416 0 17 18 0 0 4
955 206
955 220
950 220
950 243
2 12 52 0 0 12416 0 17 18 0 0 4
949 206
949 215
941 215
941 243
1 13 53 0 0 8320 0 17 18 0 0 3
943 206
932 206
932 243
2 9 54 0 0 4224 0 25 17 0 0 4
961 109
961 126
964 126
964 134
1 1 55 0 0 12416 0 20 25 0 0 4
962 62
962 67
961 67
961 73
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
