CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 120 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
143654930 0
0
6 Title:
5 Name:
0
0
0
7
7 Ground~
168 218 454 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Pulser~
4 109 471 0 10 12
0 17 18 5 19 0 0 5 5 6
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4441 0 0
0
0
6 74LS93
109 210 381 0 8 17
0 2 2 5 4 6 7 8 4
0
0 0 13040 602
6 74LS93
-21 -35 21 -27
2 U2
28 -7 42 1
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3618 0 0
0
0
6 74LS47
187 178 288 0 14 29
0 6 7 8 4 20 21 9 10 11
12 13 14 15 22
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U1
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6153 0 0
0
0
2 +V
167 193 97 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
5 DVCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
9 CA 7-Seg~
184 193 196 0 18 19
10 15 14 13 12 11 10 9 23 16
2 2 2 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7734 0 0
0
0
9 Resistor~
219 193 132 0 3 5
0 3 16 1
0
0 0 880 782
3 150
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
17
2 0 2 0 0 4096 0 3 0 0 2 3
208 411
208 423
217 423
1 1 2 0 0 4224 0 3 1 0 0 4
217 411
217 440
218 440
218 448
4 8 4 0 0 12416 0 3 3 0 0 6
190 417
190 421
175 421
175 339
190 339
190 347
3 3 5 0 0 8320 0 3 2 0 0 3
199 417
199 462
133 462
1 5 6 0 0 4224 0 4 3 0 0 4
219 325
219 339
217 339
217 347
2 6 7 0 0 4224 0 4 3 0 0 4
210 325
210 339
208 339
208 347
3 7 8 0 0 4224 0 4 3 0 0 4
201 325
201 339
199 339
199 347
4 8 4 0 0 0 0 4 3 0 0 4
192 325
192 339
190 339
190 347
7 7 9 0 0 4224 0 6 4 0 0 4
208 232
208 244
219 244
219 255
6 8 10 0 0 4224 0 6 4 0 0 4
202 232
202 250
210 250
210 255
5 9 11 0 0 4224 0 6 4 0 0 4
196 232
196 254
201 254
201 255
4 10 12 0 0 4224 0 6 4 0 0 3
190 232
190 255
192 255
3 11 13 0 0 4224 0 6 4 0 0 4
184 232
184 247
183 247
183 255
2 12 14 0 0 4224 0 6 4 0 0 4
178 232
178 256
174 256
174 255
1 13 15 0 0 4224 0 6 4 0 0 4
172 232
172 254
165 254
165 255
2 9 16 0 0 4224 0 7 6 0 0 2
193 150
193 160
1 1 3 0 0 4224 0 5 7 0 0 2
193 106
193 114
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
6227268 1079360 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
3540542 8419392 100 100 0 0
77 66 1487 276
0 447 1536 823
1487 66
77 66
1487 66
1487 276
0 0
4.53041e-315 0 4.53041e-315 0 4.53041e-315 4.53041e-315
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
